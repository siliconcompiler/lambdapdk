// //#############################################################################
// //# Function:  Positive edge-triggered static inverting D-type flop-flop with #
// //             async active low set.                                          #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_dffsqn #(
//     parameter PROP = "DEFAULT"
// ) (
//     input d,
//     input clk,
//     input nset,
//     output reg qn
// );
// 
//     always @(posedge clk or negedge nset)
//         if (!nset) qn <= 1'b0;
//         else qn <= ~d;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
module la_dffsqn (
    d,
    clk,
    nset,
    qn
);
  (* src = "generated" *)
  wire _0_;
  wire _1_;
  wire _2_;
  (* src = "generated" *)
  input clk;
  wire clk;
  (* src = "generated" *)
  input d;
  wire d;
  (* src = "generated" *)
  input nset;
  wire nset;
  (* src = "generated" *)
  output qn;
  wire qn;
  INVx2_ASAP7_75t_L _3_ (
      .A(d),
      .Y(_0_)
  );
  INVx2_ASAP7_75t_L _4_ (
      .A(_1_),
      .Y(qn)
  );
  (* src = "generated" *)
  DFFASRHQNx1_ASAP7_75t_L _5_ (
      .CLK(clk),
      .D(_0_),
      .QN(_1_),
      .RESETN(_2_),
      .SETN(nset)
  );
  TIEHIx1_ASAP7_75t_L _6_ (.H(_2_));
endmodule
