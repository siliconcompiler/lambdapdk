// //#############################################################################
// //# Function:  Positive edge-triggered static inverting D-type flop-flop with #
// //             async active low set and scan input                            #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_sdffsqn #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      si,
//     input      se,
//     input      clk,
//     input      nset,
//     output reg qn
// );
// 
//     always @(posedge clk or negedge nset)
//         if (!nset) qn <= 1'b0;
//         else qn <= se ? ~si : ~d;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_sdffsqn.v:11.1-26.10" *)
module la_sdffsqn (
    d,
    si,
    se,
    clk,
    nset,
    qn
);
  (* src = "inputs/la_sdffsqn.v:22.5-24.34" *)
  wire _0_;
  wire _1_;
  (* unused_bits = "0" *)
  wire _2_;
  (* src = "inputs/la_sdffsqn.v:17.16-17.19" *)
  input clk;
  wire clk;
  (* src = "inputs/la_sdffsqn.v:14.16-14.17" *)
  input d;
  wire d;
  (* src = "inputs/la_sdffsqn.v:18.16-18.20" *)
  input nset;
  wire nset;
  (* src = "inputs/la_sdffsqn.v:19.16-19.18" *)
  output qn;
  wire qn;
  (* src = "inputs/la_sdffsqn.v:16.16-16.18" *)
  input se;
  wire se;
  (* src = "inputs/la_sdffsqn.v:15.16-15.18" *)
  input si;
  wire si;
  MUX2_X1 _3_ (
      .A(d),
      .B(si),
      .S(se),
      .Z(_1_)
  );
  INV_X1 _4_ (
      .A (_1_),
      .ZN(_0_)
  );
  (* src = "inputs/la_sdffsqn.v:22.5-24.34" *)
  DFFR_X1 _5_ (
      .CK(clk),
      .D (_0_),
      .Q (qn),
      .QN(_2_),
      .RN(nset)
  );
endmodule
