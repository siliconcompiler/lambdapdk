// //#############################################################################
// //# Function:  Positive edge-triggered static D-type flop-flop with async     #
// //#            active low reset.                                              #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_dffrq #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      clk,
//     input      nreset,
//     output reg q
// );
// 
//     always @(posedge clk or negedge nreset)
//         if (!nreset) q <= 1'b0;
//         else q <= d;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_dffrq.v:11.1-24.10" *)
module la_dffrq (
    d,
    clk,
    nreset,
    q
);
  (* src = "inputs/la_dffrq.v:15.16-15.19" *)
  input clk;
  wire clk;
  (* src = "inputs/la_dffrq.v:14.16-14.17" *)
  input d;
  wire d;
  (* src = "inputs/la_dffrq.v:16.16-16.22" *)
  input nreset;
  wire nreset;
  (* src = "inputs/la_dffrq.v:17.16-17.17" *)
  output q;
  wire q;
  (* src = "inputs/la_dffrq.v:20.5-22.21" *)
  sky130_fd_sc_hd__dfrtp_1 _0_ (
      .CLK(clk),
      .D(d),
      .Q(q),
      .RESET_B(nreset)
  );
endmodule
