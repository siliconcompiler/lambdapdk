// //#############################################################################
// //# Function: Or-And-Inverter (oai21) Gate                                    #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_oai21 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a0,
//     input  a1,
//     input  b0,
//     output z
// );
// 
//     assign z = ~((a0 | a1) & b0);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_oai21.v:10.1-21.10" *)
module la_oai21 (
    a0,
    a1,
    b0,
    z
);
  (* src = "inputs/la_oai21.v:13.12-13.14" *)
  input a0;
  wire a0;
  (* src = "inputs/la_oai21.v:14.12-14.14" *)
  input a1;
  wire a1;
  (* src = "inputs/la_oai21.v:15.12-15.14" *)
  input b0;
  wire b0;
  (* src = "inputs/la_oai21.v:16.12-16.13" *)
  output z;
  wire z;
  sky130_fd_sc_hdll__o21ai_4 _0_ (
      .A1(a1),
      .A2(a0),
      .B1(b0),
      .Y (z)
  );
endmodule
