// //#############################################################################
// //# Function: 2-Input Inverting Mux                                           #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_muxi2 #(parameter PROP = "DEFAULT")   (
//     input  d0,
//     input  d1,
//     input  s,
//     output z
//     );
// 
//    assign z = ~((d0 & ~s) | (d1 & s));
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_muxi2(d0, d1, s, z);
  input d0;
  wire d0;
  input d1;
  wire d1;
  input s;
  wire s;
  output z;
  wire z;
  sky130_fd_sc_hd__mux2i_1 _0_ (
    .A0(d0),
    .A1(d1),
    .S(s),
    .Y(z)
  );
endmodule
