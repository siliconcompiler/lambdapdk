// //#############################################################################
// //# Function: Carry Save Adder (4:2) (aka 5:3)                                #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_csa42 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     input  b,
//     input  c,
//     input  d,
//     input  cin,
//     output sum,
//     output carry,
//     output cout
// );
// 
//     assign cout   = (a & b) | (b & c) | (a & c);
//     assign sumint = a ^ b ^ c;
//     assign sum    = cin ^ d ^ sumint;
//     assign carry  = (cin & d) | (cin & sumint) | (d & sumint);
// 
// endmodule

/* Generated by Yosys 0.38+92 (git sha1 84116c9a3, x86_64-conda-linux-gnu-cc 11.2.0 -fvisibility-inlines-hidden -fmessage-length=0 -march=nocona -mtune=haswell -ftree-vectorize -fPIC -fstack-protector-strong -fno-plt -O2 -ffunction-sections -fdebug-prefix-map=/root/conda-eda/conda-eda/workdir/conda-env/conda-bld/yosys_1708682838165/work=/usr/local/src/conda/yosys-0.38_93_g84116c9a3 -fdebug-prefix-map=/user/projekt_pia/miniconda3/envs/sc=/usr/local/src/conda-prefix -fPIC -Os -fno-merge-constants) */

module la_csa42(a, b, c, d, cin, sum, carry, cout);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  input a;
  wire a;
  input b;
  wire b;
  input c;
  wire c;
  output carry;
  wire carry;
  input cin;
  wire cin;
  output cout;
  wire cout;
  input d;
  wire d;
  output sum;
  wire sum;
  sky130_fd_sc_hdll__xnor3_1 _06_ (
    .A(b),
    .B(a),
    .C(c),
    .X(_05_)
  );
  sky130_fd_sc_hdll__xor2_1 _07_ (
    .A(d),
    .B(cin),
    .X(_00_)
  );
  sky130_fd_sc_hdll__xnor2_1 _08_ (
    .A(_05_),
    .B(_00_),
    .Y(sum)
  );
  sky130_fd_sc_hdll__nand2_6 _09_ (
    .A(d),
    .B(cin),
    .Y(_01_)
  );
  sky130_fd_sc_hdll__nor2_1 _10_ (
    .A(d),
    .B(cin),
    .Y(_02_)
  );
  sky130_fd_sc_hdll__a21oi_1 _11_ (
    .A1(_05_),
    .A2(_01_),
    .B1(_02_),
    .Y(carry)
  );
  sky130_fd_sc_hdll__nor2_1 _12_ (
    .A(b),
    .B(a),
    .Y(_03_)
  );
  sky130_fd_sc_hdll__a21oi_1 _13_ (
    .A1(b),
    .A2(a),
    .B1(c),
    .Y(_04_)
  );
  sky130_fd_sc_hdll__nor2_1 _14_ (
    .A(_03_),
    .B(_04_),
    .Y(cout)
  );
endmodule
