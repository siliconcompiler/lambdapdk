// //#############################################################################
// //# Function:  D-type active-low transparent latch                            #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_latnq #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      clk,
//     output reg q
// );
// 
//     always @(clk or d) if (~clk) q <= d;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
module la_latnq (
    d,
    clk,
    q
);
  (* src = "generated" *)
  input clk;
  wire clk;
  (* src = "generated" *)
  input d;
  wire d;
  (* src = "generated" *)
  output q;
  wire q;
  (* module_not_derived = 32'b00000000000000000000000000000001 *) (* src = "generated" *)
  DLL_X1 _0_ (
      .D (d),
      .GN(clk),
      .Q (q)
  );
endmodule
