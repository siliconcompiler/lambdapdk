// //#############################################################################
// //# Function: Or-And (oa22) Gate                                              #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_oa22 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a0,
//     input  a1,
//     input  b0,
//     input  b1,
//     output z
// );
// 
//     assign z = (a0 | a1) & (b0 | b1);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
module la_oa22 (
    a0,
    a1,
    b0,
    b1,
    z
);
  wire _0_;
  wire _1_;
  (* src = "generated" *)
  input a0;
  wire a0;
  (* src = "generated" *)
  input a1;
  wire a1;
  (* src = "generated" *)
  input b0;
  wire b0;
  (* src = "generated" *)
  input b1;
  wire b1;
  (* src = "generated" *)
  output z;
  wire z;
  sg13g2_nor2_2 _2_ (
      .A(a1),
      .B(a0),
      .Y(_0_)
  );
  sg13g2_nor2_2 _3_ (
      .A(b1),
      .B(b0),
      .Y(_1_)
  );
  sg13g2_nor2_2 _4_ (
      .A(_0_),
      .B(_1_),
      .Y(z)
  );
endmodule
