VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS

MACRO sky130_fd_sc_hdll__a2bb2o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a2bb2o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.945 0.995 1.325 1.615 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.495 0.995 1.730 1.375 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 3.365 0.765 3.625 1.655 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 2.895 1.040 3.155 1.655 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.785 0.975 1.015 ;
        RECT 0.005 0.105 3.975 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.345 2.465 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.515 2.235 0.895 2.635 ;
        RECT 2.130 2.370 2.385 2.465 ;
        RECT 1.155 2.200 2.385 2.370 ;
        RECT 2.605 2.255 2.945 2.425 ;
        RECT 1.155 1.975 1.375 2.200 ;
        RECT 0.515 1.805 1.375 1.975 ;
        RECT 2.130 2.065 2.385 2.200 ;
        RECT 0.515 0.995 0.685 1.805 ;
        RECT 1.690 1.715 1.860 1.905 ;
        RECT 2.130 1.895 2.600 2.065 ;
        RECT 1.690 1.545 2.210 1.715 ;
        RECT 2.040 0.825 2.210 1.545 ;
        RECT 1.265 0.655 2.210 0.825 ;
        RECT 2.380 0.870 2.600 1.895 ;
        RECT 2.775 2.005 2.945 2.255 ;
        RECT 3.155 2.175 3.415 2.635 ;
        RECT 3.635 2.005 3.815 2.465 ;
        RECT 2.775 1.835 3.815 2.005 ;
        RECT 2.380 0.700 2.855 0.870 ;
        RECT 0.515 0.085 0.995 0.530 ;
        RECT 1.265 0.255 1.435 0.655 ;
        RECT 1.670 0.085 2.390 0.485 ;
        RECT 2.685 0.255 2.855 0.700 ;
        RECT 3.490 0.085 3.940 0.595 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a2bb2o_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__a2bb2o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a2bb2o_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 1.445 0.995 1.815 1.615 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 1.985 0.995 2.335 1.375 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 4.080 0.765 4.455 1.655 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 3.300 1.050 3.760 1.655 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.015 0.785 1.460 1.015 ;
        RECT 0.015 0.105 4.390 0.785 ;
        RECT 0.125 -0.085 0.295 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.498000 ;
    PORT
      LAYER li1 ;
        RECT 0.525 1.525 0.830 2.465 ;
        RECT 0.525 0.810 0.745 1.525 ;
        RECT 0.525 0.255 0.830 0.810 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.185 1.445 0.355 2.635 ;
        RECT 1.000 2.235 1.380 2.635 ;
        RECT 2.700 2.370 2.870 2.465 ;
        RECT 1.640 2.200 2.870 2.370 ;
        RECT 3.125 2.255 3.455 2.425 ;
        RECT 1.640 1.975 1.860 2.200 ;
        RECT 1.000 1.805 1.860 1.975 ;
        RECT 2.640 2.065 2.870 2.200 ;
        RECT 1.000 1.325 1.220 1.805 ;
        RECT 2.175 1.715 2.345 1.905 ;
        RECT 2.640 1.895 3.100 2.065 ;
        RECT 2.175 1.545 2.710 1.715 ;
        RECT 0.915 0.995 1.220 1.325 ;
        RECT 0.185 0.085 0.355 0.930 ;
        RECT 2.540 0.825 2.710 1.545 ;
        RECT 1.765 0.655 2.710 0.825 ;
        RECT 2.880 0.870 3.100 1.895 ;
        RECT 3.285 2.005 3.455 2.255 ;
        RECT 3.675 2.175 3.925 2.635 ;
        RECT 4.145 2.005 4.315 2.465 ;
        RECT 3.285 1.835 4.315 2.005 ;
        RECT 2.880 0.700 3.280 0.870 ;
        RECT 1.000 0.085 1.480 0.530 ;
        RECT 1.765 0.255 1.935 0.655 ;
        RECT 2.155 0.085 2.890 0.485 ;
        RECT 3.110 0.255 3.280 0.700 ;
        RECT 3.905 0.085 4.355 0.595 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a2bb2o_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__a2bb2o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a2bb2o_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.820 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 3.775 1.445 5.465 1.615 ;
        RECT 3.775 1.325 4.005 1.445 ;
        RECT 3.615 1.075 4.005 1.325 ;
        RECT 5.085 1.075 5.465 1.445 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 4.205 1.075 4.915 1.275 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.445 1.835 1.615 ;
        RECT 0.085 1.075 0.625 1.445 ;
        RECT 1.665 1.245 1.835 1.445 ;
        RECT 1.665 1.075 2.095 1.245 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.855 1.075 1.445 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.820 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 7.615 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.010 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.820 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.028500 ;
    PORT
      LAYER li1 ;
        RECT 5.825 1.955 6.075 2.465 ;
        RECT 6.765 1.955 7.015 2.465 ;
        RECT 5.825 1.785 7.015 1.955 ;
        RECT 6.765 1.655 7.015 1.785 ;
        RECT 6.765 1.415 7.675 1.655 ;
        RECT 7.310 0.905 7.675 1.415 ;
        RECT 5.735 0.725 7.675 0.905 ;
        RECT 5.735 0.275 6.115 0.725 ;
        RECT 6.675 0.275 7.055 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.820 2.805 ;
        RECT 0.135 1.955 0.385 2.465 ;
        RECT 0.605 2.125 0.855 2.635 ;
        RECT 1.075 1.955 1.325 2.465 ;
        RECT 1.545 2.125 1.795 2.635 ;
        RECT 2.015 2.295 3.205 2.465 ;
        RECT 2.015 1.955 2.265 2.295 ;
        RECT 2.955 2.135 3.205 2.295 ;
        RECT 3.475 2.135 3.725 2.635 ;
        RECT 3.945 2.295 5.135 2.465 ;
        RECT 3.945 2.135 4.195 2.295 ;
        RECT 0.135 1.785 2.265 1.955 ;
        RECT 2.055 1.455 2.265 1.785 ;
        RECT 2.485 1.965 2.735 2.125 ;
        RECT 4.415 1.965 4.665 2.125 ;
        RECT 2.485 1.415 2.870 1.965 ;
        RECT 3.435 1.785 4.665 1.965 ;
        RECT 4.885 1.785 5.135 2.295 ;
        RECT 5.355 1.795 5.605 2.635 ;
        RECT 6.295 2.165 6.545 2.635 ;
        RECT 7.235 1.825 7.485 2.635 ;
        RECT 3.435 1.665 3.605 1.785 ;
        RECT 3.255 1.495 3.605 1.665 ;
        RECT 2.485 0.905 2.695 1.415 ;
        RECT 3.255 1.245 3.445 1.495 ;
        RECT 2.865 1.075 3.445 1.245 ;
        RECT 5.635 1.245 6.010 1.615 ;
        RECT 5.635 1.075 7.090 1.245 ;
        RECT 3.255 0.905 3.445 1.075 ;
        RECT 0.175 0.085 0.345 0.895 ;
        RECT 0.515 0.475 0.815 0.905 ;
        RECT 0.985 0.735 2.775 0.905 ;
        RECT 0.985 0.645 1.370 0.735 ;
        RECT 0.515 0.255 1.835 0.475 ;
        RECT 2.055 0.085 2.225 0.555 ;
        RECT 2.395 0.255 2.775 0.735 ;
        RECT 3.255 0.725 5.175 0.905 ;
        RECT 2.995 0.085 3.685 0.555 ;
        RECT 3.855 0.255 4.235 0.725 ;
        RECT 4.455 0.085 4.625 0.555 ;
        RECT 4.795 0.255 5.175 0.725 ;
        RECT 5.395 0.085 5.565 0.895 ;
        RECT 6.335 0.085 6.505 0.555 ;
        RECT 7.275 0.085 7.445 0.555 ;
        RECT 0.000 -0.085 7.820 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 2.700 1.445 2.870 1.615 ;
        RECT 5.730 1.445 5.900 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
      LAYER met1 ;
        RECT 2.640 1.600 2.980 1.645 ;
        RECT 5.670 1.600 5.960 1.645 ;
        RECT 2.640 1.460 5.960 1.600 ;
        RECT 2.640 1.415 2.980 1.460 ;
        RECT 5.670 1.415 5.960 1.460 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a2bb2o_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__a2bb2oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a2bb2oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.150 0.995 0.520 1.615 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.775 1.010 1.340 1.275 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.885 0.995 3.225 1.615 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.385 0.995 2.615 1.615 ;
        RECT 2.445 0.425 2.615 0.995 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.475 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.530000 ;
    PORT
      LAYER li1 ;
        RECT 1.520 1.955 1.885 2.465 ;
        RECT 1.520 1.785 2.155 1.955 ;
        RECT 1.985 0.825 2.155 1.785 ;
        RECT 1.985 0.255 2.275 0.825 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.095 1.805 0.425 2.635 ;
        RECT 0.925 1.615 1.305 2.465 ;
        RECT 2.055 2.235 2.495 2.465 ;
        RECT 2.325 1.955 2.495 2.235 ;
        RECT 2.665 2.135 2.915 2.635 ;
        RECT 3.135 1.955 3.390 2.465 ;
        RECT 2.325 1.785 3.390 1.955 ;
        RECT 0.925 1.445 1.815 1.615 ;
        RECT 1.645 0.830 1.815 1.445 ;
        RECT 0.095 0.085 0.425 0.825 ;
        RECT 0.645 0.660 1.815 0.830 ;
        RECT 0.645 0.255 0.815 0.660 ;
        RECT 1.045 0.085 1.715 0.490 ;
        RECT 3.005 0.085 3.385 0.825 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a2bb2oi_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__a2bb2oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a2bb2oi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 3.475 1.075 4.470 1.275 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 4.720 1.075 5.435 1.275 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.110 1.445 2.095 1.615 ;
        RECT 0.110 1.075 0.640 1.445 ;
        RECT 1.715 1.075 2.095 1.445 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.855 1.075 1.445 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.755 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.325 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.738500 ;
    PORT
      LAYER li1 ;
        RECT 2.445 0.905 2.775 2.125 ;
        RECT 0.985 0.725 2.775 0.905 ;
        RECT 0.985 0.645 1.365 0.725 ;
        RECT 2.395 0.255 2.775 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.135 1.955 0.385 2.465 ;
        RECT 0.605 2.135 0.855 2.635 ;
        RECT 1.075 1.955 1.325 2.465 ;
        RECT 1.545 2.135 1.795 2.635 ;
        RECT 2.015 2.295 3.205 2.465 ;
        RECT 2.015 1.955 2.265 2.295 ;
        RECT 0.135 1.785 2.265 1.955 ;
        RECT 2.955 1.795 3.205 2.295 ;
        RECT 3.475 1.965 3.725 2.465 ;
        RECT 3.945 2.135 4.195 2.635 ;
        RECT 4.415 2.295 5.605 2.465 ;
        RECT 4.415 1.965 4.665 2.295 ;
        RECT 3.475 1.785 4.665 1.965 ;
        RECT 4.885 1.615 5.135 2.125 ;
        RECT 3.115 1.445 5.135 1.615 ;
        RECT 5.355 1.455 5.605 2.295 ;
        RECT 3.115 1.325 3.285 1.445 ;
        RECT 2.995 0.995 3.285 1.325 ;
        RECT 3.115 0.905 3.285 0.995 ;
        RECT 0.175 0.085 0.345 0.895 ;
        RECT 0.515 0.475 0.815 0.895 ;
        RECT 3.115 0.725 5.175 0.905 ;
        RECT 0.515 0.255 1.835 0.475 ;
        RECT 2.055 0.085 2.225 0.555 ;
        RECT 2.995 0.085 3.685 0.555 ;
        RECT 3.855 0.255 4.235 0.725 ;
        RECT 4.455 0.085 4.625 0.555 ;
        RECT 4.795 0.255 5.175 0.725 ;
        RECT 5.395 0.085 5.565 0.905 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a2bb2oi_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__a2bb2oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a2bb2oi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.580 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 6.545 1.075 8.070 1.275 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 8.440 1.075 9.965 1.275 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 1.535 1.445 3.975 1.615 ;
        RECT 1.535 1.285 1.705 1.445 ;
        RECT 0.100 1.075 1.705 1.285 ;
        RECT 3.595 1.075 3.975 1.445 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 1.875 1.075 3.425 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.580 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 10.435 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.770 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.580 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.477000 ;
    PORT
      LAYER li1 ;
        RECT 4.365 1.615 4.615 2.125 ;
        RECT 5.245 1.615 5.515 2.125 ;
        RECT 4.145 1.415 5.515 1.615 ;
        RECT 4.145 0.905 4.365 1.415 ;
        RECT 1.925 0.725 5.595 0.905 ;
        RECT 1.925 0.645 3.295 0.725 ;
        RECT 4.275 0.275 4.655 0.725 ;
        RECT 5.215 0.275 5.595 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.580 2.805 ;
        RECT 0.085 1.625 0.425 2.465 ;
        RECT 0.645 1.795 0.855 2.635 ;
        RECT 1.075 1.965 1.315 2.465 ;
        RECT 1.545 2.135 1.795 2.635 ;
        RECT 2.015 1.965 2.265 2.465 ;
        RECT 2.485 2.135 2.735 2.635 ;
        RECT 2.955 1.965 3.205 2.465 ;
        RECT 3.425 2.135 3.675 2.635 ;
        RECT 3.895 2.295 6.065 2.465 ;
        RECT 3.895 1.965 4.145 2.295 ;
        RECT 1.075 1.795 4.145 1.965 ;
        RECT 4.835 1.795 5.075 2.295 ;
        RECT 1.075 1.625 1.315 1.795 ;
        RECT 0.085 1.455 1.315 1.625 ;
        RECT 5.685 1.455 6.065 2.295 ;
        RECT 6.255 1.625 6.585 2.465 ;
        RECT 6.805 1.795 7.015 2.635 ;
        RECT 7.240 1.625 7.480 2.465 ;
        RECT 7.705 1.795 7.955 2.635 ;
        RECT 8.175 2.295 10.310 2.465 ;
        RECT 8.175 1.625 8.425 2.295 ;
        RECT 6.255 1.455 8.425 1.625 ;
        RECT 8.645 1.625 8.895 2.125 ;
        RECT 9.115 1.795 9.365 2.295 ;
        RECT 9.585 1.625 9.835 2.125 ;
        RECT 10.060 1.795 10.310 2.295 ;
        RECT 8.645 1.455 10.460 1.625 ;
        RECT 4.535 1.075 6.325 1.245 ;
        RECT 6.155 0.905 6.325 1.075 ;
        RECT 10.135 0.905 10.460 1.455 ;
        RECT 0.175 0.085 0.345 0.895 ;
        RECT 0.515 0.725 1.755 0.905 ;
        RECT 6.155 0.735 10.460 0.905 ;
        RECT 0.515 0.255 0.895 0.725 ;
        RECT 1.115 0.085 1.285 0.555 ;
        RECT 1.455 0.475 1.755 0.725 ;
        RECT 6.675 0.725 9.875 0.735 ;
        RECT 1.455 0.255 3.715 0.475 ;
        RECT 3.935 0.085 4.105 0.555 ;
        RECT 4.875 0.085 5.045 0.555 ;
        RECT 5.815 0.085 6.505 0.555 ;
        RECT 6.675 0.255 7.055 0.725 ;
        RECT 7.275 0.085 7.445 0.555 ;
        RECT 7.615 0.255 7.995 0.725 ;
        RECT 8.215 0.085 8.385 0.555 ;
        RECT 8.555 0.255 8.935 0.725 ;
        RECT 9.155 0.085 9.325 0.555 ;
        RECT 9.495 0.255 9.875 0.725 ;
        RECT 10.095 0.085 10.265 0.555 ;
        RECT 0.000 -0.085 10.580 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a2bb2oi_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__a21bo_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a21bo_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.900 0.995 2.275 1.615 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.445 0.995 2.705 1.615 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.325 0.335 1.665 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.628750 ;
    PORT
      LAYER li1 ;
        RECT 3.715 0.265 3.995 2.455 ;
    END
  END X
  OBS
      LAYER pwell ;
        RECT 0.950 0.785 4.090 1.015 ;
        RECT 0.345 0.105 4.090 0.785 ;
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.105 2.045 0.345 2.435 ;
        RECT 0.515 2.225 0.915 2.635 ;
        RECT 0.105 1.845 0.965 2.045 ;
        RECT 0.515 1.165 0.965 1.845 ;
        RECT 1.135 1.345 1.465 2.455 ;
        RECT 1.685 1.985 1.865 2.455 ;
        RECT 2.035 2.155 2.415 2.635 ;
        RECT 2.640 1.985 2.810 2.455 ;
        RECT 1.685 1.785 2.810 1.985 ;
        RECT 3.075 1.495 3.360 2.635 ;
        RECT 0.515 0.265 0.795 1.165 ;
        RECT 1.135 1.045 1.730 1.345 ;
        RECT 1.045 0.085 1.290 0.865 ;
        RECT 1.460 0.815 1.730 1.045 ;
        RECT 3.285 0.815 3.545 1.325 ;
        RECT 1.460 0.625 3.545 0.815 ;
        RECT 1.460 0.265 1.940 0.625 ;
        RECT 2.620 0.085 3.350 0.455 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21bo_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__a21bo_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a21bo_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.885 0.995 3.085 1.615 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 3.375 0.995 3.665 1.615 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.225 0.995 1.695 1.325 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.965 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.547000 ;
    PORT
      LAYER li1 ;
        RECT 0.645 2.005 0.900 2.425 ;
        RECT 0.110 1.835 0.900 2.005 ;
        RECT 0.110 0.885 0.380 1.835 ;
        RECT 0.110 0.715 0.900 0.885 ;
        RECT 0.520 0.315 0.900 0.715 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.090 2.255 0.425 2.635 ;
        RECT 1.140 2.275 1.470 2.635 ;
        RECT 2.125 2.105 2.375 2.465 ;
        RECT 1.215 1.895 2.375 2.105 ;
        RECT 1.215 1.665 1.385 1.895 ;
        RECT 0.620 1.495 1.385 1.665 ;
        RECT 1.555 1.555 2.035 1.725 ;
        RECT 0.620 1.075 0.950 1.495 ;
        RECT 1.865 1.325 2.035 1.555 ;
        RECT 2.205 1.675 2.375 1.895 ;
        RECT 2.545 2.015 2.925 2.465 ;
        RECT 3.155 2.185 3.325 2.635 ;
        RECT 3.495 2.015 3.875 2.465 ;
        RECT 2.545 1.845 3.875 2.015 ;
        RECT 2.205 1.505 2.715 1.675 ;
        RECT 1.865 0.995 2.325 1.325 ;
        RECT 1.865 0.825 2.035 0.995 ;
        RECT 0.090 0.085 0.345 0.545 ;
        RECT 1.070 0.085 1.400 0.785 ;
        RECT 1.605 0.655 2.035 0.825 ;
        RECT 2.495 0.825 2.715 1.505 ;
        RECT 2.495 0.635 2.940 0.825 ;
        RECT 2.125 0.085 2.455 0.465 ;
        RECT 3.495 0.085 3.875 0.825 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21bo_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__a21bo_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a21bo_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 4.960 1.010 5.375 1.360 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 4.565 1.595 5.860 1.765 ;
        RECT 4.565 1.275 4.790 1.595 ;
        RECT 4.345 1.010 4.790 1.275 ;
        RECT 5.630 1.290 5.860 1.595 ;
        RECT 5.630 1.055 6.220 1.290 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.470 1.010 0.850 1.625 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.050 0.105 6.435 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.029000 ;
    PORT
      LAYER li1 ;
        RECT 1.050 1.595 2.580 1.765 ;
        RECT 1.050 0.785 1.540 1.595 ;
        RECT 1.050 0.615 2.510 0.785 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.105 2.105 0.520 2.465 ;
        RECT 0.690 2.275 1.070 2.635 ;
        RECT 1.650 2.275 2.030 2.635 ;
        RECT 2.605 2.275 2.990 2.635 ;
        RECT 3.275 2.210 4.385 2.380 ;
        RECT 4.555 2.275 4.935 2.635 ;
        RECT 5.495 2.275 5.875 2.635 ;
        RECT 0.105 1.935 3.090 2.105 ;
        RECT 0.105 1.795 0.535 1.935 ;
        RECT 0.105 0.840 0.300 1.795 ;
        RECT 2.920 1.525 3.090 1.935 ;
        RECT 3.275 1.695 3.445 2.210 ;
        RECT 4.205 2.105 4.385 2.210 ;
        RECT 4.205 1.935 6.345 2.105 ;
        RECT 2.920 1.355 3.525 1.525 ;
        RECT 1.710 1.185 2.750 1.325 ;
        RECT 1.710 0.995 3.030 1.185 ;
        RECT 3.215 0.995 3.525 1.355 ;
        RECT 0.105 0.255 0.510 0.840 ;
        RECT 2.860 0.785 3.030 0.995 ;
        RECT 3.745 0.840 3.915 1.805 ;
        RECT 4.205 1.445 4.385 1.935 ;
        RECT 6.090 1.460 6.345 1.935 ;
        RECT 3.745 0.785 5.385 0.840 ;
        RECT 2.860 0.670 5.385 0.785 ;
        RECT 2.860 0.615 3.915 0.670 ;
        RECT 0.680 0.085 1.070 0.445 ;
        RECT 1.650 0.085 2.030 0.445 ;
        RECT 2.735 0.085 3.505 0.445 ;
        RECT 3.745 0.255 3.915 0.615 ;
        RECT 4.175 0.085 4.505 0.445 ;
        RECT 5.105 0.405 5.385 0.670 ;
        RECT 6.065 0.085 6.345 0.885 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21bo_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__a21boi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a21boi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.985 0.375 2.240 1.345 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.650 0.995 3.125 1.345 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.975 0.335 1.665 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.885 0.785 3.165 1.015 ;
        RECT 0.295 0.105 3.165 0.785 ;
        RECT 0.295 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.676000 ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.345 1.525 2.455 ;
        RECT 1.065 1.045 1.780 1.345 ;
        RECT 1.440 0.265 1.780 1.045 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.095 2.005 0.355 2.435 ;
        RECT 0.525 2.175 0.895 2.635 ;
        RECT 0.095 1.835 0.855 2.005 ;
        RECT 0.515 0.715 0.855 1.835 ;
        RECT 1.745 1.725 1.935 2.455 ;
        RECT 2.105 1.905 2.485 2.635 ;
        RECT 2.835 1.725 3.005 2.455 ;
        RECT 1.745 1.525 3.005 1.725 ;
        RECT 0.365 0.265 0.855 0.715 ;
        RECT 1.025 0.085 1.255 0.865 ;
        RECT 2.715 0.085 3.075 0.815 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21boi_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__a21boi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a21boi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.855 0.995 3.565 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.300 1.495 4.085 1.675 ;
        RECT 2.300 1.245 2.675 1.495 ;
        RECT 2.295 1.075 2.675 1.245 ;
        RECT 3.735 0.995 4.085 1.495 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.120 0.765 0.425 1.805 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.800 0.785 4.430 1.015 ;
        RECT 0.175 0.105 4.430 0.785 ;
        RECT 0.175 0.085 0.320 0.105 ;
        RECT 0.150 -0.085 0.320 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.712500 ;
    PORT
      LAYER li1 ;
        RECT 1.525 0.785 1.865 2.115 ;
        RECT 1.525 0.615 3.360 0.785 ;
        RECT 1.525 0.255 1.870 0.615 ;
        RECT 2.980 0.255 3.360 0.615 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.095 2.080 0.425 2.635 ;
        RECT 1.100 2.285 2.415 2.465 ;
        RECT 0.645 1.285 0.825 2.265 ;
        RECT 1.100 1.795 1.350 2.285 ;
        RECT 2.035 2.025 2.415 2.285 ;
        RECT 2.635 2.195 2.805 2.635 ;
        RECT 3.110 2.105 3.280 2.465 ;
        RECT 3.460 2.275 3.840 2.635 ;
        RECT 4.060 2.105 4.320 2.465 ;
        RECT 3.110 2.025 4.320 2.105 ;
        RECT 2.035 1.855 4.320 2.025 ;
        RECT 0.645 1.070 1.355 1.285 ;
        RECT 0.645 0.530 0.825 1.070 ;
        RECT 0.265 0.360 0.825 0.530 ;
        RECT 1.085 0.085 1.325 0.885 ;
        RECT 2.140 0.085 2.470 0.445 ;
        RECT 3.990 0.085 4.330 0.785 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21boi_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__a21boi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a21boi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 3.865 1.065 5.440 1.310 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 3.300 1.480 7.120 1.705 ;
        RECT 3.300 1.065 3.695 1.480 ;
        RECT 5.725 1.075 7.120 1.480 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.075 0.670 1.615 ;
        RECT 0.450 0.995 0.670 1.075 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 7.350 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.490500 ;
    PORT
      LAYER li1 ;
        RECT 1.680 1.705 2.945 2.035 ;
        RECT 1.680 1.585 3.130 1.705 ;
        RECT 2.820 0.895 3.130 1.585 ;
        RECT 2.820 0.865 5.385 0.895 ;
        RECT 1.375 0.695 5.385 0.865 ;
        RECT 1.375 0.615 2.525 0.695 ;
        RECT 3.555 0.675 5.385 0.695 ;
        RECT 1.375 0.370 1.565 0.615 ;
        RECT 2.335 0.255 2.525 0.615 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.360 2.805 ;
        RECT 0.095 2.005 0.425 2.465 ;
        RECT 0.645 2.175 0.905 2.635 ;
        RECT 1.180 2.215 3.365 2.465 ;
        RECT 3.535 2.275 3.915 2.635 ;
        RECT 4.495 2.275 4.875 2.635 ;
        RECT 0.095 1.785 1.010 2.005 ;
        RECT 1.180 1.795 1.425 2.215 ;
        RECT 2.055 2.205 3.365 2.215 ;
        RECT 3.165 2.105 3.365 2.205 ;
        RECT 5.095 2.105 5.285 2.465 ;
        RECT 5.455 2.275 5.835 2.635 ;
        RECT 6.050 2.105 6.235 2.465 ;
        RECT 6.415 2.275 6.795 2.635 ;
        RECT 6.990 2.105 7.240 2.465 ;
        RECT 3.165 1.875 7.240 2.105 ;
        RECT 0.840 1.345 1.010 1.785 ;
        RECT 0.840 1.035 2.620 1.345 ;
        RECT 0.840 0.795 1.155 1.035 ;
        RECT 0.090 0.615 1.155 0.795 ;
        RECT 5.605 0.735 6.825 0.905 ;
        RECT 0.090 0.255 0.445 0.615 ;
        RECT 0.770 0.085 1.155 0.445 ;
        RECT 1.785 0.085 2.165 0.445 ;
        RECT 2.745 0.085 3.385 0.525 ;
        RECT 5.605 0.505 5.865 0.735 ;
        RECT 3.565 0.255 5.865 0.505 ;
        RECT 6.085 0.085 6.275 0.565 ;
        RECT 6.445 0.255 6.825 0.735 ;
        RECT 7.000 0.085 7.240 0.885 ;
        RECT 0.000 -0.085 7.360 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21boi_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__a21o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a21o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.780 1.015 2.215 1.325 ;
        RECT 1.985 0.375 2.215 1.015 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.410 0.995 2.660 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.015 1.610 1.325 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.015 0.105 2.955 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.265 0.355 2.455 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.525 1.905 0.915 2.635 ;
        RECT 1.095 1.725 1.365 2.455 ;
        RECT 0.545 1.505 1.365 1.725 ;
        RECT 1.595 1.745 1.825 2.455 ;
        RECT 2.005 1.925 2.385 2.635 ;
        RECT 2.605 1.745 2.865 2.455 ;
        RECT 1.595 1.505 2.865 1.745 ;
        RECT 0.545 0.835 0.885 1.505 ;
        RECT 0.545 0.635 1.815 0.835 ;
        RECT 0.665 0.085 1.335 0.455 ;
        RECT 1.515 0.265 1.815 0.635 ;
        RECT 2.575 0.085 2.865 0.815 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21o_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__a21o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a21o_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.410 0.365 2.730 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 3.160 0.750 3.535 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.865 0.995 2.240 1.410 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.615 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.629500 ;
    PORT
      LAYER li1 ;
        RECT 0.545 0.255 0.825 2.465 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.095 1.665 0.375 2.635 ;
        RECT 1.055 2.220 1.485 2.635 ;
        RECT 1.675 1.920 2.040 2.465 ;
        RECT 0.995 1.690 2.040 1.920 ;
        RECT 2.260 1.935 2.485 2.465 ;
        RECT 2.705 2.125 3.035 2.635 ;
        RECT 3.255 1.935 3.475 2.465 ;
        RECT 0.995 0.825 1.430 1.690 ;
        RECT 2.260 1.670 3.475 1.935 ;
        RECT 0.995 0.655 2.240 0.825 ;
        RECT 0.175 0.085 0.345 0.555 ;
        RECT 1.275 0.085 1.655 0.445 ;
        RECT 2.050 0.255 2.240 0.655 ;
        RECT 3.155 0.085 3.535 0.565 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21o_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__a21o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a21o_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 4.340 1.010 4.965 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 3.945 1.510 5.435 1.680 ;
        RECT 3.945 1.275 4.170 1.510 ;
        RECT 3.725 1.010 4.170 1.275 ;
        RECT 5.135 1.290 5.435 1.510 ;
        RECT 5.135 1.055 5.600 1.290 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.500 0.995 2.905 1.525 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.815 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.029000 ;
    PORT
      LAYER li1 ;
        RECT 0.675 1.755 0.845 2.185 ;
        RECT 1.635 1.755 1.885 2.185 ;
        RECT 0.145 1.585 1.885 1.755 ;
        RECT 0.145 0.785 0.680 1.585 ;
        RECT 0.145 0.615 1.885 0.785 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.115 1.935 0.445 2.635 ;
        RECT 1.025 1.935 1.405 2.635 ;
        RECT 2.065 1.515 2.315 2.635 ;
        RECT 2.655 2.295 3.765 2.465 ;
        RECT 2.655 1.695 2.825 2.295 ;
        RECT 0.850 0.995 2.300 1.325 ;
        RECT 2.130 0.785 2.300 0.995 ;
        RECT 3.125 0.840 3.295 2.125 ;
        RECT 3.585 2.020 3.765 2.295 ;
        RECT 3.935 2.275 4.315 2.635 ;
        RECT 4.535 2.020 4.705 2.465 ;
        RECT 4.875 2.275 5.255 2.635 ;
        RECT 5.530 2.020 5.860 2.395 ;
        RECT 3.585 1.850 5.860 2.020 ;
        RECT 3.585 1.445 3.765 1.850 ;
        RECT 5.605 1.460 5.860 1.850 ;
        RECT 3.125 0.785 4.765 0.840 ;
        RECT 2.130 0.670 4.765 0.785 ;
        RECT 2.130 0.615 3.295 0.670 ;
        RECT 0.105 0.085 0.445 0.445 ;
        RECT 1.025 0.085 1.405 0.445 ;
        RECT 2.110 0.085 2.885 0.445 ;
        RECT 3.125 0.255 3.295 0.615 ;
        RECT 3.555 0.085 3.885 0.445 ;
        RECT 4.485 0.405 4.765 0.670 ;
        RECT 5.445 0.085 5.725 0.885 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21o_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__a21o_6
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a21o_6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.900 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.865 1.055 1.535 1.290 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.525 1.460 1.875 1.630 ;
        RECT 0.525 1.290 0.695 1.460 ;
        RECT 0.095 1.055 0.695 1.290 ;
        RECT 1.705 1.290 1.875 1.460 ;
        RECT 1.705 1.055 2.045 1.290 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.865 1.055 3.195 1.615 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.900 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.115 0.105 6.645 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.090 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.900 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.396500 ;
    PORT
      LAYER li1 ;
        RECT 3.935 1.615 4.205 2.465 ;
        RECT 4.875 1.615 5.145 2.465 ;
        RECT 5.815 1.615 6.085 2.465 ;
        RECT 3.935 1.445 6.085 1.615 ;
        RECT 5.625 0.865 5.875 1.445 ;
        RECT 3.905 0.695 6.115 0.865 ;
        RECT 3.905 0.255 4.235 0.695 ;
        RECT 4.845 0.255 5.175 0.695 ;
        RECT 5.785 0.255 6.115 0.695 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.900 2.805 ;
        RECT 0.095 1.970 0.425 2.465 ;
        RECT 0.595 2.140 0.865 2.635 ;
        RECT 1.035 1.970 1.365 2.465 ;
        RECT 1.535 2.140 1.805 2.635 ;
        RECT 1.975 2.295 3.245 2.465 ;
        RECT 1.975 1.970 2.275 2.295 ;
        RECT 0.095 1.800 2.275 1.970 ;
        RECT 0.095 1.460 0.355 1.800 ;
        RECT 2.045 1.460 2.275 1.800 ;
        RECT 2.445 1.790 2.745 2.125 ;
        RECT 2.445 0.885 2.695 1.790 ;
        RECT 2.915 1.785 3.245 2.295 ;
        RECT 3.485 1.495 3.735 2.635 ;
        RECT 4.375 1.785 4.705 2.635 ;
        RECT 5.315 1.785 5.645 2.635 ;
        RECT 6.265 1.445 6.595 2.635 ;
        RECT 3.565 1.035 5.455 1.275 ;
        RECT 3.565 0.885 3.735 1.035 ;
        RECT 0.205 0.085 0.535 0.885 ;
        RECT 1.035 0.675 3.735 0.885 ;
        RECT 1.035 0.275 1.365 0.675 ;
        RECT 1.945 0.085 2.275 0.505 ;
        RECT 2.445 0.255 2.745 0.675 ;
        RECT 2.915 0.085 3.735 0.505 ;
        RECT 4.405 0.085 4.675 0.525 ;
        RECT 5.345 0.085 5.615 0.525 ;
        RECT 6.285 0.085 6.535 0.905 ;
        RECT 0.000 -0.085 6.900 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21o_6

#--------EOF---------

MACRO sky130_fd_sc_hdll__a21o_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a21o_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.820 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.865 1.055 1.535 1.290 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.525 1.460 1.875 1.630 ;
        RECT 0.525 1.290 0.695 1.460 ;
        RECT 0.095 1.055 0.695 1.290 ;
        RECT 1.705 1.290 1.875 1.460 ;
        RECT 1.705 1.055 2.045 1.290 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.865 1.055 3.195 1.615 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.820 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.115 0.105 7.585 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.010 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.820 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.862000 ;
    PORT
      LAYER li1 ;
        RECT 3.935 1.615 4.205 2.465 ;
        RECT 4.875 1.615 5.145 2.465 ;
        RECT 5.815 1.615 6.085 2.465 ;
        RECT 6.755 1.615 7.025 2.465 ;
        RECT 3.935 1.445 7.025 1.615 ;
        RECT 6.545 0.865 6.795 1.445 ;
        RECT 3.905 0.695 7.055 0.865 ;
        RECT 3.905 0.255 4.235 0.695 ;
        RECT 4.845 0.255 5.175 0.695 ;
        RECT 5.785 0.255 6.115 0.695 ;
        RECT 6.725 0.255 7.055 0.695 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.820 2.805 ;
        RECT 0.095 1.970 0.425 2.465 ;
        RECT 0.595 2.140 0.865 2.635 ;
        RECT 1.035 1.970 1.365 2.465 ;
        RECT 1.535 2.140 1.805 2.635 ;
        RECT 1.975 2.295 3.245 2.465 ;
        RECT 1.975 1.970 2.275 2.295 ;
        RECT 0.095 1.800 2.275 1.970 ;
        RECT 0.095 1.460 0.355 1.800 ;
        RECT 2.045 1.460 2.275 1.800 ;
        RECT 2.445 1.790 2.745 2.125 ;
        RECT 2.445 0.885 2.695 1.790 ;
        RECT 2.915 1.785 3.245 2.295 ;
        RECT 3.485 1.495 3.735 2.635 ;
        RECT 4.375 1.785 4.705 2.635 ;
        RECT 5.315 1.785 5.645 2.635 ;
        RECT 6.255 1.785 6.585 2.635 ;
        RECT 7.215 1.445 7.525 2.635 ;
        RECT 3.565 1.035 6.135 1.275 ;
        RECT 3.565 0.885 3.735 1.035 ;
        RECT 0.205 0.085 0.535 0.885 ;
        RECT 1.035 0.675 3.735 0.885 ;
        RECT 1.035 0.275 1.365 0.675 ;
        RECT 1.945 0.085 2.275 0.505 ;
        RECT 2.445 0.255 2.745 0.675 ;
        RECT 2.915 0.085 3.735 0.505 ;
        RECT 4.405 0.085 4.675 0.525 ;
        RECT 5.345 0.085 5.615 0.525 ;
        RECT 6.285 0.085 6.555 0.525 ;
        RECT 7.225 0.085 7.475 0.905 ;
        RECT 0.000 -0.085 7.820 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21o_8

#--------EOF---------

MACRO sky130_fd_sc_hdll__a21oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a21oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.900 0.995 1.295 1.325 ;
        RECT 1.065 0.375 1.295 0.995 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.525 0.995 1.820 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.675 0.335 1.325 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.020 0.105 1.985 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.489500 ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.685 0.370 2.455 ;
        RECT 0.095 1.495 0.730 1.685 ;
        RECT 0.505 0.825 0.730 1.495 ;
        RECT 0.505 0.645 0.885 0.825 ;
        RECT 0.660 0.265 0.885 0.645 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.540 2.025 0.920 2.455 ;
        RECT 1.140 2.195 1.335 2.635 ;
        RECT 1.515 2.025 1.895 2.455 ;
        RECT 0.540 1.855 1.895 2.025 ;
        RECT 0.900 1.525 1.895 1.855 ;
        RECT 0.110 0.085 0.440 0.475 ;
        RECT 1.595 0.085 1.895 0.815 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21oi_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__a21oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a21oi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.895 0.995 1.575 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.145 1.495 2.130 1.675 ;
        RECT 0.145 1.035 0.695 1.495 ;
        RECT 1.755 1.075 2.130 1.495 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 3.035 0.995 3.535 1.625 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.515 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.745000 ;
    PORT
      LAYER li1 ;
        RECT 2.515 1.330 2.865 2.115 ;
        RECT 2.410 0.785 2.865 1.330 ;
        RECT 1.005 0.615 2.865 0.785 ;
        RECT 1.005 0.255 1.400 0.615 ;
        RECT 2.545 0.255 2.865 0.615 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.110 2.105 0.370 2.465 ;
        RECT 0.540 2.275 0.920 2.635 ;
        RECT 1.150 2.105 1.320 2.465 ;
        RECT 1.625 2.195 1.795 2.635 ;
        RECT 2.015 2.285 3.390 2.465 ;
        RECT 0.110 2.025 1.320 2.105 ;
        RECT 2.015 2.025 2.345 2.285 ;
        RECT 0.110 1.855 2.345 2.025 ;
        RECT 3.085 1.795 3.390 2.285 ;
        RECT 0.100 0.085 0.395 0.865 ;
        RECT 1.910 0.085 2.290 0.445 ;
        RECT 3.095 0.085 3.425 0.825 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21oi_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__a21oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a21oi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 2.815 1.065 4.400 1.310 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 2.250 1.480 6.070 1.705 ;
        RECT 2.250 1.065 2.645 1.480 ;
        RECT 4.675 1.075 6.070 1.480 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.035 1.580 1.415 ;
        RECT 0.090 0.995 0.400 1.035 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 6.315 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.523000 ;
    PORT
      LAYER li1 ;
        RECT 0.630 1.705 1.895 2.035 ;
        RECT 0.630 1.585 2.080 1.705 ;
        RECT 1.750 0.895 2.080 1.585 ;
        RECT 1.750 0.865 4.305 0.895 ;
        RECT 0.645 0.695 4.305 0.865 ;
        RECT 0.645 0.615 1.795 0.695 ;
        RECT 2.475 0.675 4.305 0.695 ;
        RECT 0.645 0.370 0.835 0.615 ;
        RECT 1.605 0.255 1.795 0.615 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.180 2.215 2.315 2.465 ;
        RECT 2.485 2.275 2.865 2.635 ;
        RECT 0.180 1.795 0.375 2.215 ;
        RECT 1.005 2.205 2.315 2.215 ;
        RECT 2.115 2.105 2.315 2.205 ;
        RECT 3.085 2.105 3.275 2.465 ;
        RECT 3.445 2.275 3.825 2.635 ;
        RECT 4.045 2.105 4.235 2.465 ;
        RECT 4.405 2.275 4.785 2.635 ;
        RECT 5.005 2.105 5.185 2.465 ;
        RECT 5.365 2.275 5.745 2.635 ;
        RECT 5.965 2.105 6.225 2.465 ;
        RECT 2.115 1.875 6.225 2.105 ;
        RECT 0.090 0.085 0.425 0.805 ;
        RECT 4.525 0.735 5.745 0.905 ;
        RECT 1.005 0.085 1.385 0.445 ;
        RECT 1.985 0.085 2.315 0.525 ;
        RECT 4.525 0.505 4.785 0.735 ;
        RECT 2.485 0.255 4.785 0.505 ;
        RECT 5.005 0.085 5.195 0.565 ;
        RECT 5.365 0.255 5.745 0.735 ;
        RECT 5.965 0.085 6.225 0.885 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21oi_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__a22o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a22o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.525 1.065 2.085 1.285 ;
        RECT 1.525 0.675 1.745 1.065 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.275 0.980 2.625 1.285 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.815 1.075 1.285 1.285 ;
        RECT 1.065 0.675 1.285 1.075 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.625 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.615 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.670000 ;
    PORT
      LAYER li1 ;
        RECT 3.275 1.785 3.535 2.465 ;
        RECT 3.365 0.585 3.535 1.785 ;
        RECT 3.275 0.255 3.535 0.585 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.090 2.245 0.425 2.465 ;
        RECT 1.540 2.255 1.895 2.635 ;
        RECT 0.090 1.715 0.345 2.245 ;
        RECT 2.065 2.085 2.395 2.465 ;
        RECT 0.565 1.885 2.395 2.085 ;
        RECT 2.585 1.935 2.915 2.635 ;
        RECT 0.090 1.495 3.035 1.715 ;
        RECT 0.090 0.085 0.595 0.850 ;
        RECT 2.865 0.785 3.035 1.495 ;
        RECT 2.110 0.615 3.035 0.785 ;
        RECT 2.110 0.465 2.280 0.615 ;
        RECT 0.870 0.255 2.280 0.465 ;
        RECT 2.585 0.085 2.915 0.445 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a22o_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__a22o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a22o_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.525 1.075 1.940 1.285 ;
        RECT 1.525 0.675 1.820 1.075 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.160 1.075 2.615 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.815 1.075 1.340 1.285 ;
        RECT 1.065 0.675 1.340 1.075 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 0.625 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.095 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.498000 ;
    PORT
      LAYER li1 ;
        RECT 3.150 1.785 3.560 2.465 ;
        RECT 3.240 0.585 3.560 1.785 ;
        RECT 3.150 0.255 3.560 0.585 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.095 2.295 1.365 2.465 ;
        RECT 0.095 1.625 0.425 2.295 ;
        RECT 1.035 2.255 1.365 2.295 ;
        RECT 1.555 2.215 1.910 2.635 ;
        RECT 0.645 2.035 0.875 2.125 ;
        RECT 2.130 2.035 2.380 2.465 ;
        RECT 0.645 1.795 2.380 2.035 ;
        RECT 2.600 1.875 2.930 2.635 ;
        RECT 0.095 1.455 3.015 1.625 ;
        RECT 2.845 0.905 3.015 1.455 ;
        RECT 3.755 1.445 3.925 2.635 ;
        RECT 0.095 0.085 0.595 0.850 ;
        RECT 2.125 0.735 3.015 0.905 ;
        RECT 2.125 0.505 2.295 0.735 ;
        RECT 0.870 0.255 2.295 0.505 ;
        RECT 2.505 0.085 2.885 0.565 ;
        RECT 3.755 0.085 3.925 0.985 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a22o_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__a22o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a22o_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.900 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 5.350 1.075 5.895 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 4.750 1.445 6.285 1.615 ;
        RECT 4.750 1.075 5.130 1.445 ;
        RECT 6.115 1.275 6.285 1.445 ;
        RECT 6.115 1.075 6.815 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 3.375 1.075 4.030 1.275 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.620 1.445 4.580 1.615 ;
        RECT 2.620 1.075 3.205 1.445 ;
        RECT 4.200 1.075 4.580 1.445 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.900 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.070 0.105 6.840 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.090 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.900 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.028500 ;
    PORT
      LAYER li1 ;
        RECT 0.690 1.615 0.940 2.465 ;
        RECT 1.630 1.615 1.880 2.465 ;
        RECT 0.085 1.445 1.880 1.615 ;
        RECT 0.085 0.905 0.370 1.445 ;
        RECT 0.085 0.725 1.920 0.905 ;
        RECT 0.600 0.265 0.980 0.725 ;
        RECT 1.540 0.255 1.920 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.900 2.805 ;
        RECT 0.220 1.825 0.470 2.635 ;
        RECT 1.160 1.795 1.410 2.635 ;
        RECT 2.100 2.125 2.350 2.635 ;
        RECT 2.620 2.295 4.830 2.465 ;
        RECT 2.620 2.125 2.870 2.295 ;
        RECT 3.560 2.125 3.810 2.295 ;
        RECT 3.090 1.955 3.340 2.125 ;
        RECT 4.030 1.955 4.280 2.125 ;
        RECT 2.100 1.785 4.280 1.955 ;
        RECT 4.500 1.955 4.830 2.295 ;
        RECT 5.050 2.125 5.300 2.635 ;
        RECT 5.520 1.955 5.770 2.465 ;
        RECT 5.990 2.125 6.240 2.635 ;
        RECT 6.505 1.955 6.710 2.465 ;
        RECT 4.500 1.785 6.710 1.955 ;
        RECT 2.100 1.275 2.430 1.785 ;
        RECT 6.505 1.455 6.710 1.785 ;
        RECT 0.540 1.075 2.430 1.275 ;
        RECT 2.140 0.905 2.430 1.075 ;
        RECT 2.140 0.735 5.810 0.905 ;
        RECT 3.420 0.645 3.905 0.735 ;
        RECT 5.385 0.645 5.810 0.735 ;
        RECT 0.260 0.085 0.430 0.555 ;
        RECT 1.200 0.085 1.370 0.555 ;
        RECT 2.140 0.085 2.830 0.555 ;
        RECT 3.000 0.255 4.320 0.475 ;
        RECT 4.585 0.085 4.755 0.555 ;
        RECT 6.030 0.475 6.280 0.895 ;
        RECT 4.960 0.255 6.280 0.475 ;
        RECT 6.500 0.085 6.670 0.895 ;
        RECT 0.000 -0.085 6.900 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a22o_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__a22oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a22oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.525 1.055 2.085 1.275 ;
        RECT 1.525 0.675 1.735 1.055 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.265 0.995 2.625 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.815 1.075 1.315 1.275 ;
        RECT 1.065 0.675 1.315 1.075 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.765 0.625 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.955 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.917000 ;
    PORT
      LAYER li1 ;
        RECT 0.095 2.295 1.375 2.465 ;
        RECT 0.095 1.615 0.425 2.295 ;
        RECT 1.035 2.195 1.375 2.295 ;
        RECT 0.095 1.445 3.135 1.615 ;
        RECT 2.795 0.825 3.135 1.445 ;
        RECT 2.095 0.655 3.135 0.825 ;
        RECT 2.095 0.505 2.275 0.655 ;
        RECT 0.870 0.255 2.275 0.505 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 1.555 2.255 1.910 2.635 ;
        RECT 0.645 1.980 0.815 2.115 ;
        RECT 2.105 1.980 2.275 2.165 ;
        RECT 0.645 1.785 2.275 1.980 ;
        RECT 2.560 1.855 2.825 2.635 ;
        RECT 0.095 0.085 0.595 0.595 ;
        RECT 2.505 0.085 2.835 0.485 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a22oi_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__a22oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a22oi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.645 1.075 3.535 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 3.770 1.075 4.620 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 1.030 1.075 1.745 1.275 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.150 1.075 0.830 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.895 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.278500 ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.655 0.345 2.465 ;
        RECT 0.985 1.655 1.365 2.125 ;
        RECT 1.925 1.655 2.360 2.125 ;
        RECT 0.095 1.485 2.360 1.655 ;
        RECT 1.930 0.845 2.360 1.485 ;
        RECT 1.455 0.675 3.295 0.845 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.060 2.805 ;
        RECT 0.515 2.295 2.825 2.465 ;
        RECT 0.515 1.825 0.815 2.295 ;
        RECT 1.585 1.825 1.755 2.295 ;
        RECT 2.575 1.655 2.825 2.295 ;
        RECT 3.045 1.825 3.215 2.635 ;
        RECT 3.385 1.655 3.865 2.465 ;
        RECT 4.085 1.825 4.255 2.635 ;
        RECT 4.425 1.655 4.805 2.465 ;
        RECT 2.575 1.485 4.805 1.655 ;
        RECT 0.095 0.680 1.285 0.850 ;
        RECT 0.095 0.255 0.345 0.680 ;
        RECT 0.515 0.085 0.895 0.510 ;
        RECT 1.115 0.505 1.285 0.680 ;
        RECT 3.615 0.680 4.875 0.850 ;
        RECT 3.615 0.505 3.785 0.680 ;
        RECT 1.115 0.255 2.305 0.505 ;
        RECT 2.495 0.255 3.785 0.505 ;
        RECT 3.980 0.085 4.360 0.510 ;
        RECT 4.555 0.255 4.875 0.680 ;
        RECT 0.000 -0.085 5.060 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a22oi_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__a22oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a22oi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.740 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 4.675 1.075 6.285 1.285 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 6.510 1.075 8.535 1.285 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 2.865 1.075 4.440 1.275 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 2.095 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.740 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 8.555 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.930 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.740 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.024500 ;
    PORT
      LAYER li1 ;
        RECT 0.645 1.625 0.855 2.125 ;
        RECT 1.545 1.625 1.795 2.125 ;
        RECT 2.485 1.625 2.735 2.125 ;
        RECT 3.425 1.625 3.675 2.125 ;
        RECT 0.645 1.445 3.675 1.625 ;
        RECT 2.395 0.885 2.695 1.445 ;
        RECT 2.395 0.645 6.115 0.885 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.740 2.805 ;
        RECT 0.090 2.295 4.665 2.465 ;
        RECT 0.090 1.455 0.425 2.295 ;
        RECT 1.075 1.795 1.325 2.295 ;
        RECT 2.015 1.795 2.265 2.295 ;
        RECT 2.955 1.795 3.205 2.295 ;
        RECT 3.895 1.625 4.665 2.295 ;
        RECT 4.885 1.795 5.135 2.635 ;
        RECT 5.355 1.625 5.605 2.465 ;
        RECT 5.825 1.795 6.075 2.635 ;
        RECT 6.295 1.625 6.545 2.465 ;
        RECT 6.765 1.795 7.015 2.635 ;
        RECT 7.235 1.625 7.485 2.465 ;
        RECT 7.705 1.795 7.955 2.635 ;
        RECT 8.175 1.625 8.425 2.465 ;
        RECT 3.895 1.455 8.425 1.625 ;
        RECT 0.095 0.725 2.225 0.905 ;
        RECT 0.095 0.255 0.425 0.725 ;
        RECT 0.645 0.085 0.815 0.555 ;
        RECT 0.985 0.255 1.365 0.725 ;
        RECT 1.585 0.085 1.755 0.555 ;
        RECT 1.925 0.475 2.225 0.725 ;
        RECT 6.335 0.725 8.465 0.905 ;
        RECT 6.335 0.475 6.585 0.725 ;
        RECT 1.925 0.255 4.185 0.475 ;
        RECT 4.375 0.255 6.585 0.475 ;
        RECT 6.805 0.085 6.975 0.555 ;
        RECT 7.145 0.255 7.525 0.725 ;
        RECT 7.745 0.085 7.915 0.555 ;
        RECT 8.085 0.255 8.465 0.725 ;
        RECT 0.000 -0.085 8.740 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a22oi_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__a31o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a31o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.985 0.995 2.275 1.655 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.515 0.995 1.815 1.655 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.075 1.325 1.340 1.655 ;
        RECT 0.985 0.995 1.340 1.325 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.445 0.995 2.745 1.655 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.175 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.447250 ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.575 0.425 2.425 ;
        RECT 0.095 0.810 0.285 1.575 ;
        RECT 0.095 0.300 0.425 0.810 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.645 1.495 0.895 2.635 ;
        RECT 1.085 1.995 1.385 2.415 ;
        RECT 1.665 2.165 1.995 2.635 ;
        RECT 2.275 1.995 2.525 2.415 ;
        RECT 1.085 1.825 2.525 1.995 ;
        RECT 2.755 1.825 3.085 2.425 ;
        RECT 0.455 0.995 0.815 1.325 ;
        RECT 0.645 0.825 0.815 0.995 ;
        RECT 2.915 0.825 3.085 1.825 ;
        RECT 0.645 0.655 3.085 0.825 ;
        RECT 0.605 0.085 0.935 0.485 ;
        RECT 2.125 0.315 2.505 0.655 ;
        RECT 2.725 0.085 3.055 0.485 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a31o_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__a31o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a31o_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.385 0.415 2.615 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.905 0.400 2.155 1.325 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.030 0.995 1.545 1.325 ;
        RECT 1.030 0.760 1.370 0.995 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 3.195 0.755 3.535 1.325 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.545 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.530500 ;
    PORT
      LAYER li1 ;
        RECT 0.645 2.005 0.815 2.465 ;
        RECT 0.090 1.835 0.815 2.005 ;
        RECT 0.090 0.885 0.345 1.835 ;
        RECT 0.090 0.715 0.815 0.885 ;
        RECT 0.645 0.255 0.815 0.715 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.135 2.175 0.385 2.635 ;
        RECT 0.985 1.835 1.285 2.635 ;
        RECT 1.455 2.005 1.755 2.425 ;
        RECT 2.015 2.175 2.345 2.635 ;
        RECT 2.585 2.005 2.895 2.425 ;
        RECT 1.455 1.835 2.895 2.005 ;
        RECT 3.175 1.665 3.345 2.465 ;
        RECT 0.515 1.495 3.345 1.665 ;
        RECT 0.515 1.245 0.685 1.495 ;
        RECT 0.515 1.075 0.845 1.245 ;
        RECT 0.090 0.085 0.425 0.465 ;
        RECT 1.005 0.085 1.385 0.465 ;
        RECT 2.785 0.255 2.955 1.495 ;
        RECT 3.175 0.085 3.465 0.565 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a31o_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__a31o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a31o_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.900 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 1.455 1.075 1.855 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.775 0.905 1.255 1.275 ;
        RECT 2.185 1.075 2.565 1.275 ;
        RECT 2.185 0.905 2.370 1.075 ;
        RECT 0.775 0.735 2.370 0.905 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.145 1.445 3.155 1.615 ;
        RECT 0.145 1.075 0.525 1.445 ;
        RECT 2.775 1.075 3.155 1.445 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 3.925 1.075 4.455 1.285 ;
        RECT 4.215 0.745 4.455 1.075 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.900 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 6.795 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.090 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.900 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.996000 ;
    PORT
      LAYER li1 ;
        RECT 5.045 1.955 5.215 2.465 ;
        RECT 5.985 1.955 6.155 2.465 ;
        RECT 4.935 1.785 6.780 1.955 ;
        RECT 6.585 0.825 6.780 1.785 ;
        RECT 4.905 0.655 6.780 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.900 2.805 ;
        RECT 0.175 1.955 0.345 2.465 ;
        RECT 0.515 2.125 0.895 2.635 ;
        RECT 1.115 1.955 1.285 2.465 ;
        RECT 1.455 2.125 1.835 2.635 ;
        RECT 2.055 1.955 2.225 2.465 ;
        RECT 2.395 2.125 2.775 2.635 ;
        RECT 3.115 2.295 4.225 2.465 ;
        RECT 3.115 1.955 3.285 2.295 ;
        RECT 0.175 1.785 3.285 1.955 ;
        RECT 3.455 1.625 3.835 2.115 ;
        RECT 4.055 1.795 4.225 2.295 ;
        RECT 4.495 2.125 4.825 2.635 ;
        RECT 5.385 2.125 5.765 2.635 ;
        RECT 6.325 2.125 6.705 2.635 ;
        RECT 3.455 1.455 4.820 1.625 ;
        RECT 0.175 0.085 0.345 0.905 ;
        RECT 3.455 0.870 3.695 1.455 ;
        RECT 4.650 1.325 4.820 1.455 ;
        RECT 4.650 0.995 6.355 1.325 ;
        RECT 2.600 0.805 3.695 0.870 ;
        RECT 2.600 0.700 3.835 0.805 ;
        RECT 2.600 0.565 2.770 0.700 ;
        RECT 1.455 0.395 2.770 0.565 ;
        RECT 2.950 0.085 3.285 0.530 ;
        RECT 3.455 0.295 3.835 0.700 ;
        RECT 4.135 0.085 4.665 0.565 ;
        RECT 5.385 0.085 5.765 0.485 ;
        RECT 6.325 0.085 6.705 0.485 ;
        RECT 0.000 -0.085 6.900 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a31o_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__a31oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a31oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.445 1.695 1.665 ;
        RECT 1.370 0.995 1.695 1.445 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.335 1.165 1.275 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.435 1.325 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.325 0.995 2.650 1.325 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.665 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.523750 ;
    PORT
      LAYER li1 ;
        RECT 1.985 1.495 2.410 2.445 ;
        RECT 1.985 0.825 2.155 1.495 ;
        RECT 1.480 0.295 2.155 0.825 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.090 1.495 0.420 2.635 ;
        RECT 0.640 2.005 0.815 2.415 ;
        RECT 1.035 2.175 1.365 2.635 ;
        RECT 1.620 2.005 1.815 2.415 ;
        RECT 0.640 1.835 1.815 2.005 ;
        RECT 0.090 0.085 0.430 0.815 ;
        RECT 2.325 0.085 2.585 0.565 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a31oi_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__a31oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a31oi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.330 0.995 3.090 1.615 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 1.150 0.995 1.905 1.615 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.995 0.870 1.615 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 4.715 1.275 4.940 1.625 ;
        RECT 4.220 1.075 4.940 1.275 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.045 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.007000 ;
    PORT
      LAYER li1 ;
        RECT 4.155 1.615 4.485 2.115 ;
        RECT 3.330 1.445 4.485 1.615 ;
        RECT 3.330 0.845 3.645 1.445 ;
        RECT 3.330 0.825 4.955 0.845 ;
        RECT 2.545 0.655 4.955 0.825 ;
        RECT 3.605 0.255 3.775 0.655 ;
        RECT 4.575 0.295 4.955 0.655 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.060 2.805 ;
        RECT 0.175 1.955 0.345 2.465 ;
        RECT 0.515 2.125 0.895 2.635 ;
        RECT 1.115 1.955 1.285 2.465 ;
        RECT 1.455 2.125 1.835 2.635 ;
        RECT 2.055 1.955 2.225 2.465 ;
        RECT 2.560 2.125 3.280 2.635 ;
        RECT 3.685 2.295 4.875 2.465 ;
        RECT 3.685 1.955 3.855 2.295 ;
        RECT 0.175 1.785 3.855 1.955 ;
        RECT 4.705 1.795 4.875 2.295 ;
        RECT 0.095 0.655 2.305 0.825 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.455 0.295 3.375 0.465 ;
        RECT 4.025 0.085 4.405 0.465 ;
        RECT 0.000 -0.085 5.060 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a31oi_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__a31oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a31oi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.740 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 4.225 0.995 6.020 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 2.135 0.995 3.950 1.325 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.120 0.995 1.885 1.325 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 6.270 0.995 7.605 1.630 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.740 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 8.665 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.930 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.740 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.613500 ;
    PORT
      LAYER li1 ;
        RECT 6.725 1.915 8.085 2.085 ;
        RECT 7.845 0.805 8.085 1.915 ;
        RECT 4.425 0.635 8.435 0.805 ;
        RECT 7.325 0.255 7.495 0.635 ;
        RECT 8.265 0.255 8.435 0.635 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.740 2.805 ;
        RECT 0.175 1.665 0.345 2.465 ;
        RECT 0.515 1.915 0.895 2.635 ;
        RECT 1.115 1.665 1.285 2.465 ;
        RECT 1.455 1.915 1.835 2.635 ;
        RECT 2.055 1.665 2.225 2.465 ;
        RECT 2.395 1.915 2.775 2.635 ;
        RECT 2.995 1.665 3.165 2.465 ;
        RECT 3.335 1.915 3.715 2.635 ;
        RECT 3.935 1.665 4.105 2.465 ;
        RECT 4.295 1.915 4.675 2.635 ;
        RECT 4.895 1.665 5.065 2.465 ;
        RECT 5.235 2.255 5.615 2.635 ;
        RECT 5.835 2.425 6.005 2.465 ;
        RECT 5.835 2.255 8.515 2.425 ;
        RECT 5.835 1.665 6.005 2.255 ;
        RECT 0.175 1.495 6.005 1.665 ;
        RECT 8.265 1.495 8.515 2.255 ;
        RECT 0.175 0.635 4.185 0.805 ;
        RECT 0.175 0.255 0.345 0.635 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.115 0.255 1.285 0.635 ;
        RECT 1.455 0.085 1.835 0.465 ;
        RECT 2.055 0.255 2.225 0.635 ;
        RECT 2.395 0.295 6.165 0.465 ;
        RECT 6.725 0.085 7.105 0.465 ;
        RECT 7.665 0.085 8.045 0.465 ;
        RECT 0.000 -0.085 8.740 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a31oi_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__a32o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a32o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.260 0.955 2.665 1.325 ;
        RECT 2.380 0.665 2.665 0.955 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.525 0.665 1.950 1.325 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.015 0.995 1.355 1.325 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.835 0.660 3.135 1.325 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 3.790 1.325 4.030 1.615 ;
        RECT 3.430 0.995 4.030 1.325 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.975 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.554500 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.915 0.425 2.425 ;
        RECT 0.090 0.560 0.345 1.915 ;
        RECT 0.090 0.300 0.425 0.560 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.725 1.835 1.055 2.635 ;
        RECT 1.350 2.045 1.635 2.465 ;
        RECT 1.940 2.215 2.270 2.635 ;
        RECT 2.545 2.295 3.895 2.465 ;
        RECT 2.545 2.045 2.875 2.295 ;
        RECT 1.350 1.875 2.875 2.045 ;
        RECT 3.155 1.665 3.325 2.125 ;
        RECT 3.635 1.795 3.895 2.295 ;
        RECT 0.675 1.495 3.325 1.665 ;
        RECT 0.675 1.325 0.845 1.495 ;
        RECT 0.570 0.995 0.845 1.325 ;
        RECT 0.675 0.825 0.845 0.995 ;
        RECT 0.675 0.655 1.315 0.825 ;
        RECT 1.145 0.485 1.315 0.655 ;
        RECT 0.595 0.085 0.975 0.485 ;
        RECT 1.145 0.315 2.910 0.485 ;
        RECT 3.505 0.085 3.885 0.805 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a32o_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__a32o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a32o_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.875 0.415 3.145 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 3.315 0.425 3.650 1.625 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 4.165 0.995 4.505 1.630 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.245 2.670 1.615 ;
        RECT 2.235 1.075 2.670 1.245 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.065 0.745 1.630 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.485 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.748000 ;
    PORT
      LAYER li1 ;
        RECT 0.135 1.955 0.345 2.465 ;
        RECT 1.115 1.955 1.285 2.465 ;
        RECT 0.135 1.785 1.285 1.955 ;
        RECT 0.135 0.825 0.345 1.785 ;
        RECT 0.135 0.655 0.895 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.515 2.125 0.895 2.635 ;
        RECT 1.635 2.295 2.745 2.465 ;
        RECT 1.635 1.785 1.805 2.295 ;
        RECT 2.025 1.945 2.355 2.115 ;
        RECT 2.575 1.965 2.745 2.295 ;
        RECT 2.915 2.140 3.295 2.635 ;
        RECT 3.675 1.965 3.845 2.465 ;
        RECT 2.025 1.615 2.275 1.945 ;
        RECT 2.575 1.795 3.845 1.965 ;
        RECT 4.015 1.915 4.400 2.635 ;
        RECT 0.535 1.445 2.275 1.615 ;
        RECT 0.535 0.995 0.755 1.445 ;
        RECT 1.800 0.845 2.040 1.445 ;
        RECT 1.800 0.675 2.705 0.845 ;
        RECT 0.090 0.085 0.425 0.465 ;
        RECT 0.985 0.085 1.740 0.445 ;
        RECT 2.405 0.295 2.705 0.675 ;
        RECT 4.015 0.085 4.400 0.805 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a32o_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__a32o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a32o_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.280 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 4.680 1.075 5.575 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 3.635 1.075 4.430 1.325 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.410 1.075 3.405 1.295 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 6.120 1.075 7.140 1.625 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 7.440 1.295 7.635 1.635 ;
        RECT 7.440 1.075 8.170 1.295 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.280 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 8.275 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.470 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.280 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.028500 ;
    PORT
      LAYER li1 ;
        RECT 0.645 1.665 0.815 2.465 ;
        RECT 1.585 1.665 1.755 2.465 ;
        RECT 0.120 1.495 1.755 1.665 ;
        RECT 0.120 0.805 0.340 1.495 ;
        RECT 0.120 0.635 1.755 0.805 ;
        RECT 0.645 0.255 0.815 0.635 ;
        RECT 1.585 0.255 1.755 0.635 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.280 2.805 ;
        RECT 0.095 1.915 0.425 2.635 ;
        RECT 0.985 1.915 1.365 2.635 ;
        RECT 1.925 1.915 2.305 2.635 ;
        RECT 2.525 2.085 2.695 2.465 ;
        RECT 2.865 2.255 3.245 2.635 ;
        RECT 3.515 2.085 3.685 2.465 ;
        RECT 3.855 2.255 4.235 2.635 ;
        RECT 4.455 2.085 4.625 2.465 ;
        RECT 4.795 2.255 5.175 2.635 ;
        RECT 5.395 2.255 8.185 2.425 ;
        RECT 5.395 2.085 5.565 2.255 ;
        RECT 2.525 1.915 5.565 2.085 ;
        RECT 6.445 2.075 7.715 2.085 ;
        RECT 5.780 1.915 7.715 2.075 ;
        RECT 5.780 1.905 6.510 1.915 ;
        RECT 5.780 1.665 5.950 1.905 ;
        RECT 7.935 1.755 8.185 2.255 ;
        RECT 1.950 1.495 5.950 1.665 ;
        RECT 1.950 1.325 2.170 1.495 ;
        RECT 0.620 0.995 2.170 1.325 ;
        RECT 2.525 0.655 4.235 0.825 ;
        RECT 5.780 0.805 5.950 1.495 ;
        RECT 0.095 0.085 0.425 0.465 ;
        RECT 0.985 0.085 1.365 0.465 ;
        RECT 1.925 0.085 2.305 0.465 ;
        RECT 2.525 0.255 2.695 0.655 ;
        RECT 4.795 0.635 6.735 0.805 ;
        RECT 6.995 0.645 8.105 0.815 ;
        RECT 6.995 0.465 7.165 0.645 ;
        RECT 2.865 0.085 3.245 0.465 ;
        RECT 3.435 0.295 5.645 0.465 ;
        RECT 5.930 0.295 7.165 0.465 ;
        RECT 6.995 0.255 7.165 0.295 ;
        RECT 7.335 0.085 7.715 0.465 ;
        RECT 7.935 0.255 8.105 0.645 ;
        RECT 0.000 -0.085 8.280 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a32o_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__a32oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a32oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.475 0.345 1.695 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.985 0.415 2.185 1.325 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.390 1.015 2.855 1.325 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.945 0.995 1.235 1.615 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.345 1.325 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.035 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.634500 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.785 0.915 2.085 ;
        RECT 0.515 0.805 0.775 1.785 ;
        RECT 0.515 0.635 1.265 0.805 ;
        RECT 0.965 0.295 1.265 0.635 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.085 2.255 1.445 2.465 ;
        RECT 0.085 1.835 0.345 2.255 ;
        RECT 1.195 1.955 1.445 2.255 ;
        RECT 1.705 2.135 1.955 2.635 ;
        RECT 2.215 1.955 2.385 2.465 ;
        RECT 1.195 1.785 2.385 1.955 ;
        RECT 2.215 1.745 2.385 1.785 ;
        RECT 2.555 1.495 2.945 2.635 ;
        RECT 0.110 0.085 0.440 0.465 ;
        RECT 2.570 0.085 2.960 0.805 ;
        RECT 0.000 -0.085 3.235 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a32oi_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__a32oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a32oi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.375 1.075 3.255 1.625 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 3.720 1.075 4.575 1.625 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 5.025 1.075 6.320 1.625 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.075 1.795 1.285 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.145 1.285 0.325 1.625 ;
        RECT 0.145 1.075 0.875 1.285 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 6.435 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.195 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.996000 ;
    PORT
      LAYER li1 ;
        RECT 0.565 1.625 0.895 2.125 ;
        RECT 1.585 1.625 1.755 2.125 ;
        RECT 0.565 1.455 2.195 1.625 ;
        RECT 1.965 0.825 2.195 1.455 ;
        RECT 1.455 0.655 3.245 0.825 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.175 2.295 2.225 2.465 ;
        RECT 0.175 1.795 0.345 2.295 ;
        RECT 1.115 1.795 1.285 2.295 ;
        RECT 2.055 1.965 2.225 2.295 ;
        RECT 2.445 2.255 3.165 2.635 ;
        RECT 3.415 1.965 3.585 2.465 ;
        RECT 3.770 2.255 4.525 2.635 ;
        RECT 4.695 1.965 4.865 2.465 ;
        RECT 5.125 2.255 5.845 2.635 ;
        RECT 6.095 1.965 6.265 2.465 ;
        RECT 2.055 1.795 6.265 1.965 ;
        RECT 0.095 0.715 1.285 0.885 ;
        RECT 0.095 0.295 0.425 0.715 ;
        RECT 0.645 0.085 0.815 0.545 ;
        RECT 1.035 0.465 1.285 0.715 ;
        RECT 3.755 0.635 5.800 0.805 ;
        RECT 1.035 0.295 2.305 0.465 ;
        RECT 2.495 0.295 4.605 0.465 ;
        RECT 4.865 0.085 5.250 0.465 ;
        RECT 5.420 0.275 5.800 0.635 ;
        RECT 6.095 0.085 6.265 0.885 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a32oi_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__a32oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a32oi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.500 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 4.175 1.075 6.065 1.285 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 6.745 1.075 8.545 1.300 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 9.145 1.075 11.035 1.280 ;
        RECT 10.755 0.755 11.035 1.075 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 2.835 0.995 3.955 1.325 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.110 1.305 0.330 1.965 ;
        RECT 0.110 1.075 1.900 1.305 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.500 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 11.165 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 11.690 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.500 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.024500 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.745 0.895 2.085 ;
        RECT 1.455 1.745 1.835 2.085 ;
        RECT 2.175 1.745 2.775 2.085 ;
        RECT 3.335 1.745 3.715 2.085 ;
        RECT 0.515 1.575 3.715 1.745 ;
        RECT 2.175 0.990 2.615 1.575 ;
        RECT 2.395 0.805 2.615 0.990 ;
        RECT 2.395 0.635 6.165 0.805 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 11.500 2.805 ;
        RECT 0.095 2.255 4.105 2.425 ;
        RECT 3.935 1.745 4.105 2.255 ;
        RECT 4.295 1.915 4.675 2.635 ;
        RECT 4.895 1.745 5.065 2.465 ;
        RECT 5.320 1.915 6.040 2.635 ;
        RECT 6.290 1.745 6.460 2.465 ;
        RECT 6.865 1.915 7.245 2.635 ;
        RECT 7.465 1.745 7.635 2.465 ;
        RECT 7.805 1.915 8.185 2.635 ;
        RECT 8.405 1.745 8.575 2.465 ;
        RECT 9.265 1.915 9.645 2.635 ;
        RECT 9.865 1.745 10.035 2.465 ;
        RECT 10.205 1.915 10.585 2.635 ;
        RECT 10.805 1.745 10.975 2.465 ;
        RECT 3.935 1.575 10.975 1.745 ;
        RECT 0.175 0.635 2.225 0.805 ;
        RECT 6.865 0.635 10.505 0.805 ;
        RECT 0.175 0.255 0.345 0.635 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.115 0.255 1.285 0.635 ;
        RECT 2.055 0.465 2.225 0.635 ;
        RECT 1.455 0.085 1.835 0.465 ;
        RECT 2.055 0.295 4.185 0.465 ;
        RECT 4.425 0.295 8.655 0.465 ;
        RECT 8.845 0.085 9.175 0.465 ;
        RECT 9.395 0.255 9.565 0.635 ;
        RECT 9.735 0.085 10.115 0.465 ;
        RECT 10.335 0.255 10.505 0.635 ;
        RECT 10.685 0.085 11.075 0.465 ;
        RECT 0.000 -0.085 11.500 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a32oi_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__a211o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a211o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.865 0.995 2.390 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.015 0.995 1.695 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.590 0.995 3.075 1.325 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 3.305 0.995 3.585 1.325 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.665 1.015 ;
        RECT 0.135 -0.085 0.305 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.447250 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.685 0.355 2.455 ;
        RECT 0.090 0.265 0.425 1.685 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.525 1.915 0.905 2.635 ;
        RECT 1.095 2.095 1.355 2.455 ;
        RECT 1.525 2.265 2.085 2.635 ;
        RECT 2.305 2.095 2.565 2.455 ;
        RECT 1.095 1.865 2.565 2.095 ;
        RECT 3.205 1.685 3.545 2.455 ;
        RECT 0.605 1.505 3.545 1.685 ;
        RECT 0.605 0.815 0.845 1.505 ;
        RECT 0.605 0.625 3.535 0.815 ;
        RECT 0.655 0.085 1.400 0.455 ;
        RECT 2.195 0.265 2.520 0.625 ;
        RECT 2.700 0.085 3.080 0.455 ;
        RECT 3.310 0.265 3.535 0.625 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a211o_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__a211o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a211o_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.290 1.045 2.695 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.525 1.045 1.960 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.865 1.045 3.195 1.275 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 3.365 1.045 3.735 1.275 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.025 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.504500 ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.255 0.835 2.335 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.090 1.490 0.385 2.635 ;
        RECT 1.100 1.830 1.355 2.635 ;
        RECT 1.555 2.020 1.935 2.465 ;
        RECT 2.155 2.190 2.430 2.635 ;
        RECT 2.715 2.020 3.045 2.465 ;
        RECT 1.555 1.840 3.045 2.020 ;
        RECT 3.555 1.660 3.935 2.325 ;
        RECT 1.100 1.490 3.935 1.660 ;
        RECT 0.090 0.085 0.385 0.905 ;
        RECT 1.100 0.875 1.355 1.490 ;
        RECT 1.100 0.695 3.935 0.875 ;
        RECT 1.005 0.085 1.770 0.445 ;
        RECT 2.475 0.275 2.855 0.695 ;
        RECT 3.110 0.085 3.385 0.525 ;
        RECT 3.555 0.275 3.935 0.695 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a211o_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__a211o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a211o_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 5.535 1.020 5.930 1.330 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 4.945 1.510 6.445 1.700 ;
        RECT 4.945 1.020 5.325 1.510 ;
        RECT 6.125 1.320 6.445 1.510 ;
        RECT 6.125 1.020 6.875 1.320 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.875 1.445 4.625 1.700 ;
        RECT 2.875 1.325 3.105 1.445 ;
        RECT 2.790 0.985 3.105 1.325 ;
        RECT 4.245 0.985 4.625 1.445 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 3.275 0.985 4.045 1.275 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.071250 ;
    PORT
      LAYER li1 ;
        RECT 0.645 1.705 0.830 2.465 ;
        RECT 1.600 1.705 1.790 2.465 ;
        RECT 0.085 1.495 1.790 1.705 ;
        RECT 0.085 0.875 0.340 1.495 ;
        RECT 0.085 0.635 2.225 0.875 ;
        RECT 1.085 0.615 2.225 0.635 ;
        RECT 1.085 0.255 1.275 0.615 ;
        RECT 2.045 0.255 2.225 0.615 ;
    END
  END X
  OBS
      LAYER pwell ;
        RECT 0.395 0.105 7.085 1.015 ;
      LAYER li1 ;
        RECT 0.000 2.635 7.360 2.805 ;
        RECT 0.090 1.875 0.425 2.635 ;
        RECT 1.050 1.875 1.380 2.635 ;
        RECT 2.010 1.835 2.260 2.635 ;
        RECT 2.570 2.210 4.900 2.465 ;
        RECT 5.070 2.275 5.450 2.635 ;
        RECT 4.570 2.105 4.900 2.210 ;
        RECT 5.660 2.105 5.970 2.465 ;
        RECT 6.140 2.275 6.520 2.635 ;
        RECT 6.740 2.105 6.995 2.465 ;
        RECT 2.530 1.870 3.860 2.040 ;
        RECT 4.570 1.880 6.995 2.105 ;
        RECT 2.530 1.675 2.705 1.870 ;
        RECT 2.385 1.505 2.705 1.675 ;
        RECT 6.615 1.535 6.995 1.880 ;
        RECT 2.385 1.325 2.620 1.505 ;
        RECT 0.525 1.045 2.620 1.325 ;
        RECT 2.395 0.805 2.620 1.045 ;
        RECT 2.395 0.615 6.040 0.805 ;
        RECT 0.485 0.085 0.865 0.465 ;
        RECT 1.445 0.085 1.825 0.445 ;
        RECT 2.420 0.085 2.805 0.445 ;
        RECT 3.025 0.255 3.270 0.615 ;
        RECT 3.440 0.085 3.820 0.445 ;
        RECT 4.040 0.255 4.420 0.615 ;
        RECT 4.640 0.085 5.010 0.445 ;
        RECT 5.660 0.275 6.040 0.615 ;
        RECT 6.615 0.085 6.995 0.805 ;
        RECT 0.000 -0.085 7.360 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a211o_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__a211oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a211oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.995 1.280 1.325 ;
        RECT 0.605 0.265 0.905 0.995 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.765 0.435 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.500 0.995 1.795 2.455 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.980 0.995 2.265 1.615 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.610 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.870250 ;
    PORT
      LAYER li1 ;
        RECT 1.965 1.785 2.650 2.455 ;
        RECT 2.435 0.815 2.650 1.785 ;
        RECT 1.155 0.625 2.650 0.815 ;
        RECT 1.155 0.265 1.340 0.625 ;
        RECT 2.255 0.265 2.480 0.625 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.125 1.725 0.375 2.455 ;
        RECT 0.545 1.905 0.925 2.635 ;
        RECT 1.145 1.725 1.330 2.455 ;
        RECT 0.125 1.525 1.330 1.725 ;
        RECT 0.085 0.085 0.425 0.595 ;
        RECT 1.550 0.085 1.930 0.455 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a211oi_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__a211oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a211oi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.810 1.035 3.570 1.285 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 4.685 1.285 4.915 1.655 ;
        RECT 3.890 1.035 4.915 1.285 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.285 1.285 1.615 ;
        RECT 1.065 1.035 1.935 1.285 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.100 0.995 0.405 1.615 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.055 0.105 4.925 1.015 ;
        RECT 0.125 -0.085 0.295 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008500 ;
    PORT
      LAYER li1 ;
        RECT 0.575 0.855 0.895 2.115 ;
        RECT 0.575 0.655 3.395 0.855 ;
        RECT 0.575 0.255 0.885 0.655 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.060 2.805 ;
        RECT 0.145 2.285 2.415 2.455 ;
        RECT 0.145 1.785 0.405 2.285 ;
        RECT 1.175 2.255 2.415 2.285 ;
        RECT 1.175 1.785 1.365 2.255 ;
        RECT 1.535 1.655 1.915 2.075 ;
        RECT 2.135 1.835 2.415 2.255 ;
        RECT 2.635 1.835 2.865 2.635 ;
        RECT 3.095 1.655 3.365 2.465 ;
        RECT 3.595 1.835 3.825 2.635 ;
        RECT 4.055 1.655 4.325 2.465 ;
        RECT 4.555 1.835 4.785 2.635 ;
        RECT 1.535 1.455 4.325 1.655 ;
        RECT 0.145 0.085 0.395 0.815 ;
        RECT 3.625 0.635 4.835 0.855 ;
        RECT 3.625 0.475 3.795 0.635 ;
        RECT 1.055 0.085 1.435 0.475 ;
        RECT 2.015 0.085 2.395 0.475 ;
        RECT 2.585 0.265 3.795 0.475 ;
        RECT 3.975 0.085 4.355 0.455 ;
        RECT 4.585 0.265 4.835 0.635 ;
        RECT 0.000 -0.085 5.060 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a211oi_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__a211oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a211oi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.280 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 1.805 1.035 3.305 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.100 1.445 3.975 1.625 ;
        RECT 0.100 1.035 1.535 1.445 ;
        RECT 3.595 1.035 3.975 1.445 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER met1 ;
        RECT 4.225 1.600 4.515 1.645 ;
        RECT 7.280 1.600 7.570 1.645 ;
        RECT 4.225 1.460 7.570 1.600 ;
        RECT 4.225 1.415 4.515 1.460 ;
        RECT 7.280 1.415 7.570 1.460 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 6.830 1.275 7.050 1.695 ;
        RECT 5.550 1.035 7.050 1.275 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.280 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 8.155 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.470 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.280 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.985000 ;
    PORT
      LAYER li1 ;
        RECT 5.720 1.865 8.160 2.085 ;
        RECT 7.680 1.495 8.160 1.865 ;
        RECT 1.925 0.825 7.055 0.865 ;
        RECT 7.905 0.825 8.160 1.495 ;
        RECT 1.925 0.695 8.160 0.825 ;
        RECT 1.925 0.675 3.680 0.695 ;
        RECT 4.275 0.625 8.160 0.695 ;
        RECT 4.275 0.615 5.595 0.625 ;
        RECT 4.275 0.255 4.645 0.615 ;
        RECT 5.425 0.255 5.595 0.615 ;
        RECT 6.365 0.615 8.160 0.625 ;
        RECT 6.365 0.255 6.535 0.615 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.280 2.805 ;
        RECT 0.095 2.085 0.345 2.465 ;
        RECT 0.515 2.255 0.895 2.635 ;
        RECT 1.115 2.105 1.285 2.465 ;
        RECT 1.455 2.275 1.835 2.635 ;
        RECT 2.055 2.105 2.225 2.465 ;
        RECT 2.395 2.275 2.775 2.635 ;
        RECT 2.995 2.105 3.165 2.465 ;
        RECT 3.335 2.275 3.715 2.635 ;
        RECT 3.935 2.255 8.070 2.465 ;
        RECT 3.935 2.105 4.105 2.255 ;
        RECT 1.115 2.085 4.105 2.105 ;
        RECT 0.095 1.795 4.105 2.085 ;
        RECT 4.275 1.785 5.460 2.085 ;
        RECT 5.130 1.695 5.460 1.785 ;
        RECT 4.145 1.275 4.960 1.615 ;
        RECT 5.130 1.445 6.610 1.695 ;
        RECT 7.300 1.325 7.510 1.655 ;
        RECT 4.145 1.035 5.305 1.275 ;
        RECT 7.300 0.995 7.735 1.325 ;
        RECT 0.615 0.695 1.755 0.865 ;
        RECT 0.095 0.085 0.395 0.585 ;
        RECT 0.615 0.530 0.825 0.695 ;
        RECT 1.000 0.085 1.285 0.525 ;
        RECT 1.455 0.505 1.755 0.695 ;
        RECT 1.455 0.255 3.715 0.505 ;
        RECT 3.935 0.085 4.105 0.525 ;
        RECT 4.865 0.085 5.195 0.445 ;
        RECT 5.815 0.085 6.145 0.445 ;
        RECT 6.755 0.085 7.085 0.445 ;
        RECT 7.665 0.085 8.070 0.445 ;
        RECT 0.000 -0.085 8.280 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 4.285 1.445 4.455 1.615 ;
        RECT 7.340 1.445 7.510 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a211oi_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__a221oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a221oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.985 1.075 2.425 1.285 ;
        RECT 1.985 0.675 2.350 1.075 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.670 0.995 3.075 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.325 1.075 1.815 1.285 ;
        RECT 1.525 0.675 1.815 1.075 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.075 1.155 1.285 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.435 1.285 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.470 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.874500 ;
    PORT
      LAYER li1 ;
        RECT 0.175 1.625 0.345 2.465 ;
        RECT 2.300 1.625 3.535 1.665 ;
        RECT 0.175 1.495 3.535 1.625 ;
        RECT 0.175 1.455 2.450 1.495 ;
        RECT 0.170 0.735 1.335 0.905 ;
        RECT 3.255 0.825 3.535 1.495 ;
        RECT 0.170 0.255 0.345 0.735 ;
        RECT 1.165 0.505 1.335 0.735 ;
        RECT 2.580 0.655 3.535 0.825 ;
        RECT 2.580 0.505 2.780 0.655 ;
        RECT 1.165 0.255 2.780 0.505 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.515 2.295 1.835 2.465 ;
        RECT 0.515 1.795 0.815 2.295 ;
        RECT 1.455 2.255 1.835 2.295 ;
        RECT 2.025 2.215 2.355 2.635 ;
        RECT 1.115 2.045 1.340 2.125 ;
        RECT 2.575 2.045 2.825 2.465 ;
        RECT 1.115 1.835 2.825 2.045 ;
        RECT 3.045 1.875 3.375 2.635 ;
        RECT 1.115 1.795 2.175 1.835 ;
        RECT 0.515 0.085 0.895 0.565 ;
        RECT 3.030 0.085 3.360 0.485 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a221oi_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__a221oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a221oi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 4.235 1.075 4.915 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 3.735 1.445 5.270 1.615 ;
        RECT 3.735 1.075 4.065 1.445 ;
        RECT 5.100 1.275 5.270 1.445 ;
        RECT 5.100 1.075 5.885 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.360 1.075 3.015 1.275 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 1.730 1.445 3.565 1.615 ;
        RECT 1.730 1.075 2.190 1.445 ;
        RECT 3.185 1.075 3.565 1.445 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 0.420 1.615 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.825 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.979000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.905 0.905 2.125 ;
        RECT 0.605 0.865 4.795 0.905 ;
        RECT 0.525 0.725 4.795 0.865 ;
        RECT 0.525 0.305 0.905 0.725 ;
        RECT 2.435 0.645 2.835 0.725 ;
        RECT 4.415 0.645 4.795 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.090 2.295 1.375 2.465 ;
        RECT 0.090 1.795 0.435 2.295 ;
        RECT 1.125 1.955 1.375 2.295 ;
        RECT 1.605 2.295 3.775 2.465 ;
        RECT 1.605 2.125 1.855 2.295 ;
        RECT 2.545 2.125 2.795 2.295 ;
        RECT 2.075 1.955 2.325 2.125 ;
        RECT 3.015 1.955 3.265 2.125 ;
        RECT 1.125 1.785 3.265 1.955 ;
        RECT 3.525 1.955 3.775 2.295 ;
        RECT 4.035 2.125 4.285 2.635 ;
        RECT 4.505 1.955 4.755 2.465 ;
        RECT 4.975 2.125 5.225 2.635 ;
        RECT 5.490 1.955 5.695 2.465 ;
        RECT 3.525 1.785 5.695 1.955 ;
        RECT 1.125 1.495 1.375 1.785 ;
        RECT 5.490 1.455 5.695 1.785 ;
        RECT 0.105 0.085 0.355 0.895 ;
        RECT 1.125 0.085 1.815 0.555 ;
        RECT 1.985 0.255 3.305 0.475 ;
        RECT 3.570 0.085 3.740 0.555 ;
        RECT 5.015 0.475 5.265 0.905 ;
        RECT 3.945 0.255 5.265 0.475 ;
        RECT 5.485 0.085 5.655 0.905 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a221oi_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__a221oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a221oi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.580 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 7.145 1.075 8.755 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 6.585 1.445 9.135 1.615 ;
        RECT 6.585 1.075 6.965 1.445 ;
        RECT 8.965 1.275 9.135 1.445 ;
        RECT 8.965 1.075 10.400 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 4.335 0.995 5.885 1.275 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 3.945 1.445 6.410 1.615 ;
        RECT 3.945 1.325 4.165 1.445 ;
        RECT 3.765 0.995 4.165 1.325 ;
        RECT 6.065 1.075 6.410 1.445 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 1.435 1.275 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.580 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 10.530 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.770 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.580 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.893000 ;
    PORT
      LAYER li1 ;
        RECT 0.625 1.615 0.875 2.125 ;
        RECT 1.565 1.615 1.815 2.125 ;
        RECT 0.625 1.445 1.855 1.615 ;
        RECT 1.655 1.275 1.855 1.445 ;
        RECT 1.655 1.095 3.595 1.275 ;
        RECT 1.655 0.905 1.855 1.095 ;
        RECT 0.535 0.725 1.855 0.905 ;
        RECT 0.535 0.255 0.915 0.725 ;
        RECT 1.475 0.255 1.855 0.725 ;
        RECT 3.375 0.820 3.595 1.095 ;
        RECT 6.110 0.820 7.130 0.905 ;
        RECT 3.375 0.735 8.585 0.820 ;
        RECT 3.375 0.645 6.280 0.735 ;
        RECT 6.960 0.645 8.585 0.735 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.580 2.805 ;
        RECT 0.090 2.295 2.325 2.465 ;
        RECT 0.090 1.445 0.405 2.295 ;
        RECT 1.095 1.785 1.345 2.295 ;
        RECT 2.075 1.615 2.325 2.295 ;
        RECT 2.565 2.215 6.655 2.465 ;
        RECT 6.825 2.215 9.085 2.635 ;
        RECT 2.565 1.795 2.815 2.215 ;
        RECT 6.405 2.045 6.655 2.215 ;
        RECT 9.275 2.045 9.445 2.465 ;
        RECT 3.035 1.835 6.185 2.045 ;
        RECT 3.035 1.615 3.330 1.835 ;
        RECT 6.405 1.785 9.525 2.045 ;
        RECT 9.745 1.795 9.915 2.635 ;
        RECT 2.075 1.445 3.330 1.615 ;
        RECT 9.355 1.615 9.525 1.785 ;
        RECT 10.175 1.615 10.425 2.465 ;
        RECT 9.355 1.445 10.425 1.615 ;
        RECT 0.115 0.085 0.365 0.895 ;
        RECT 2.075 0.645 3.205 0.925 ;
        RECT 1.135 0.085 1.305 0.555 ;
        RECT 2.075 0.085 2.245 0.645 ;
        RECT 3.035 0.595 3.205 0.645 ;
        RECT 8.805 0.725 9.995 0.905 ;
        RECT 2.435 0.425 2.860 0.475 ;
        RECT 3.335 0.425 6.185 0.475 ;
        RECT 2.435 0.255 6.185 0.425 ;
        RECT 6.455 0.085 6.625 0.555 ;
        RECT 8.805 0.475 9.055 0.725 ;
        RECT 6.795 0.255 9.055 0.475 ;
        RECT 9.275 0.085 9.445 0.555 ;
        RECT 9.615 0.255 9.995 0.725 ;
        RECT 10.165 0.085 10.335 0.905 ;
        RECT 0.000 -0.085 10.580 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a221oi_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__a222oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a222oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.276000 ;
    PORT
      LAYER li1 ;
        RECT 2.905 1.000 3.305 1.330 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.276000 ;
    PORT
      LAYER li1 ;
        RECT 3.475 1.000 3.995 1.330 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.276000 ;
    PORT
      LAYER li1 ;
        RECT 2.415 1.000 2.735 1.330 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.276000 ;
    PORT
      LAYER li1 ;
        RECT 1.885 1.000 2.245 1.330 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.276000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.000 0.595 1.315 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.276000 ;
    PORT
      LAYER li1 ;
        RECT 0.765 1.000 1.235 1.315 ;
    END
  END C2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.105 1.005 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.981600 ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.795 0.345 2.295 ;
        RECT 0.095 1.485 1.655 1.795 ;
        RECT 1.405 0.815 1.655 1.485 ;
        RECT 0.095 0.645 2.975 0.815 ;
        RECT 0.095 0.255 0.425 0.645 ;
        RECT 2.410 0.295 2.975 0.645 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.565 2.295 2.465 2.465 ;
        RECT 0.565 2.055 0.895 2.295 ;
        RECT 2.170 2.135 2.465 2.295 ;
        RECT 2.685 1.830 2.935 2.250 ;
        RECT 3.155 1.905 3.485 2.635 ;
        RECT 1.825 1.735 2.935 1.830 ;
        RECT 3.765 1.735 4.025 2.250 ;
        RECT 1.825 1.500 4.025 1.735 ;
        RECT 0.925 0.085 1.705 0.465 ;
        RECT 3.555 0.085 3.965 0.815 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a222oi_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__and2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.100 1.325 0.455 1.685 ;
        RECT 0.100 1.075 0.665 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.885 1.075 1.235 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.040 0.925 2.085 1.015 ;
        RECT 0.005 0.245 2.085 0.925 ;
        RECT 0.145 0.105 2.085 0.245 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.757250 ;
    PORT
      LAYER li1 ;
        RECT 1.730 1.915 2.155 2.465 ;
        RECT 1.860 0.545 2.155 1.915 ;
        RECT 1.525 0.255 2.155 0.545 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.125 1.965 0.405 2.635 ;
        RECT 0.625 1.745 0.925 2.295 ;
        RECT 1.095 1.915 1.425 2.635 ;
        RECT 0.625 1.575 1.575 1.745 ;
        RECT 1.405 1.325 1.575 1.575 ;
        RECT 1.405 0.995 1.660 1.325 ;
        RECT 1.405 0.905 1.575 0.995 ;
        RECT 0.125 0.715 1.575 0.905 ;
        RECT 0.125 0.355 0.455 0.715 ;
        RECT 1.105 0.085 1.355 0.545 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and2_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__and2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.325 0.350 1.765 ;
        RECT 0.095 1.075 0.715 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.885 1.075 1.265 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.085 0.925 2.735 1.015 ;
        RECT 0.005 0.245 2.735 0.925 ;
        RECT 0.145 0.105 2.735 0.245 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.728500 ;
    PORT
      LAYER li1 ;
        RECT 1.745 1.915 2.205 2.465 ;
        RECT 1.935 0.545 2.205 1.915 ;
        RECT 1.595 0.255 2.205 0.545 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.115 1.965 0.395 2.635 ;
        RECT 0.615 1.745 0.915 2.295 ;
        RECT 1.165 1.915 1.505 2.635 ;
        RECT 0.615 1.575 1.605 1.745 ;
        RECT 1.435 1.325 1.605 1.575 ;
        RECT 2.375 1.495 2.665 2.635 ;
        RECT 1.435 0.995 1.765 1.325 ;
        RECT 1.435 0.905 1.605 0.995 ;
        RECT 0.115 0.715 1.605 0.905 ;
        RECT 0.115 0.355 0.445 0.715 ;
        RECT 1.175 0.085 1.425 0.545 ;
        RECT 2.375 0.085 2.665 0.885 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and2_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__and2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.995 0.435 1.615 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.995 1.080 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.490 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.061500 ;
    PORT
      LAYER li1 ;
        RECT 1.680 1.760 1.870 2.465 ;
        RECT 2.640 1.765 2.830 2.465 ;
        RECT 2.640 1.760 3.570 1.765 ;
        RECT 1.680 1.535 3.570 1.760 ;
        RECT 3.290 0.845 3.570 1.535 ;
        RECT 1.680 0.615 3.570 0.845 ;
        RECT 1.680 0.515 1.870 0.615 ;
        RECT 2.640 0.255 2.830 0.615 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.095 1.880 0.425 2.635 ;
        RECT 0.655 1.750 0.835 2.465 ;
        RECT 1.090 1.935 1.420 2.635 ;
        RECT 2.040 1.935 2.420 2.635 ;
        RECT 3.000 1.935 3.380 2.635 ;
        RECT 0.655 1.580 1.460 1.750 ;
        RECT 1.250 1.355 1.460 1.580 ;
        RECT 1.250 1.020 2.935 1.355 ;
        RECT 1.250 0.805 1.460 1.020 ;
        RECT 0.095 0.615 1.460 0.805 ;
        RECT 0.095 0.255 0.425 0.615 ;
        RECT 1.055 0.085 1.385 0.445 ;
        RECT 2.040 0.085 2.420 0.445 ;
        RECT 3.000 0.085 3.380 0.445 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and2_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__and2_6
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and2_6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.865 0.995 1.535 1.295 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.435 1.465 1.885 1.635 ;
        RECT 0.435 1.325 0.615 1.465 ;
        RECT 0.085 0.995 0.615 1.325 ;
        RECT 1.705 1.325 1.885 1.465 ;
        RECT 1.705 0.995 1.965 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.235 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.396500 ;
    PORT
      LAYER li1 ;
        RECT 2.475 1.615 2.745 2.465 ;
        RECT 3.415 1.615 3.685 2.465 ;
        RECT 4.355 1.615 4.625 2.465 ;
        RECT 2.475 1.445 4.975 1.615 ;
        RECT 4.475 0.885 4.975 1.445 ;
        RECT 2.475 0.715 4.975 0.885 ;
        RECT 2.475 0.255 2.745 0.715 ;
        RECT 3.415 0.255 3.685 0.715 ;
        RECT 4.355 0.255 4.625 0.715 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.095 1.805 0.395 2.635 ;
        RECT 0.565 1.975 0.865 2.465 ;
        RECT 1.035 2.145 1.365 2.635 ;
        RECT 1.535 1.975 1.805 2.465 ;
        RECT 1.975 2.160 2.305 2.635 ;
        RECT 0.565 1.805 2.305 1.975 ;
        RECT 2.135 1.265 2.305 1.805 ;
        RECT 2.915 1.785 3.245 2.635 ;
        RECT 3.855 1.785 4.185 2.635 ;
        RECT 4.795 1.785 5.125 2.635 ;
        RECT 2.135 1.055 4.305 1.265 ;
        RECT 2.135 0.825 2.305 1.055 ;
        RECT 0.095 0.085 0.425 0.825 ;
        RECT 1.015 0.655 2.305 0.825 ;
        RECT 1.015 0.255 1.345 0.655 ;
        RECT 1.940 0.085 2.270 0.485 ;
        RECT 2.915 0.085 3.245 0.545 ;
        RECT 3.855 0.085 4.185 0.545 ;
        RECT 4.795 0.085 5.125 0.545 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and2_6

#--------EOF---------

MACRO sky130_fd_sc_hdll__and2_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and2_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.865 0.995 1.535 1.295 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.435 1.465 1.885 1.635 ;
        RECT 0.435 1.325 0.615 1.465 ;
        RECT 0.085 0.995 0.615 1.325 ;
        RECT 1.705 1.325 1.885 1.465 ;
        RECT 1.705 0.995 1.965 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 6.175 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.862000 ;
    PORT
      LAYER li1 ;
        RECT 2.475 1.615 2.745 2.465 ;
        RECT 3.415 1.615 3.685 2.465 ;
        RECT 4.355 1.615 4.625 2.465 ;
        RECT 5.295 1.615 5.565 2.465 ;
        RECT 2.475 1.445 5.915 1.615 ;
        RECT 5.495 0.885 5.915 1.445 ;
        RECT 2.475 0.715 5.915 0.885 ;
        RECT 2.475 0.255 2.745 0.715 ;
        RECT 3.415 0.255 3.685 0.715 ;
        RECT 4.355 0.255 4.625 0.715 ;
        RECT 5.295 0.255 5.565 0.715 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.095 1.805 0.395 2.635 ;
        RECT 0.565 1.975 0.865 2.465 ;
        RECT 1.035 2.145 1.365 2.635 ;
        RECT 1.535 1.975 1.805 2.465 ;
        RECT 1.975 2.160 2.305 2.635 ;
        RECT 0.565 1.805 2.305 1.975 ;
        RECT 2.135 1.265 2.305 1.805 ;
        RECT 2.915 1.785 3.245 2.635 ;
        RECT 3.855 1.785 4.185 2.635 ;
        RECT 4.795 1.785 5.125 2.635 ;
        RECT 5.735 1.785 6.065 2.635 ;
        RECT 2.135 1.055 5.325 1.265 ;
        RECT 2.135 0.825 2.305 1.055 ;
        RECT 0.095 0.085 0.425 0.825 ;
        RECT 1.015 0.655 2.305 0.825 ;
        RECT 1.015 0.255 1.345 0.655 ;
        RECT 1.940 0.085 2.270 0.485 ;
        RECT 2.915 0.085 3.245 0.545 ;
        RECT 3.855 0.085 4.185 0.545 ;
        RECT 4.795 0.085 5.125 0.545 ;
        RECT 5.735 0.085 6.065 0.545 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and2_8

#--------EOF---------

MACRO sky130_fd_sc_hdll__and2b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and2b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.765 0.445 1.615 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.630 1.645 2.275 1.955 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.025 0.785 3.045 1.015 ;
        RECT 0.005 0.105 3.045 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.505000 ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.580 3.080 2.365 ;
        RECT 2.770 0.775 3.080 1.580 ;
        RECT 2.705 0.255 3.080 0.775 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.175 2.015 0.345 2.445 ;
        RECT 0.515 2.185 0.895 2.635 ;
        RECT 0.175 1.785 0.900 2.015 ;
        RECT 0.665 1.135 0.900 1.785 ;
        RECT 1.070 1.475 1.405 2.420 ;
        RECT 1.635 2.165 2.275 2.635 ;
        RECT 1.070 1.325 2.080 1.475 ;
        RECT 1.070 1.305 2.505 1.325 ;
        RECT 0.665 0.805 1.250 1.135 ;
        RECT 1.420 0.945 2.505 1.305 ;
        RECT 0.665 0.655 0.885 0.805 ;
        RECT 0.090 0.085 0.425 0.590 ;
        RECT 0.645 0.280 0.885 0.655 ;
        RECT 1.420 0.610 1.640 0.945 ;
        RECT 1.215 0.415 1.640 0.610 ;
        RECT 1.215 0.270 1.385 0.415 ;
        RECT 2.000 0.085 2.445 0.580 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and2b_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__and2b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and2b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.765 0.450 1.615 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.655 1.645 2.400 1.955 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.050 0.785 3.675 1.015 ;
        RECT 0.005 0.105 3.675 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.762000 ;
    PORT
      LAYER li1 ;
        RECT 2.575 1.580 3.090 2.365 ;
        RECT 2.755 0.775 3.090 1.580 ;
        RECT 2.695 0.255 3.090 0.775 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.175 2.015 0.345 2.445 ;
        RECT 0.515 2.185 0.895 2.635 ;
        RECT 0.175 1.785 0.905 2.015 ;
        RECT 0.670 1.135 0.905 1.785 ;
        RECT 1.095 1.475 1.430 2.420 ;
        RECT 1.660 2.165 2.395 2.635 ;
        RECT 3.325 1.680 3.595 2.635 ;
        RECT 1.095 1.325 2.105 1.475 ;
        RECT 1.095 1.305 2.535 1.325 ;
        RECT 0.670 0.805 1.275 1.135 ;
        RECT 1.445 0.945 2.535 1.305 ;
        RECT 0.670 0.655 0.885 0.805 ;
        RECT 0.095 0.085 0.425 0.590 ;
        RECT 0.645 0.280 0.885 0.655 ;
        RECT 1.445 0.610 1.665 0.945 ;
        RECT 1.215 0.415 1.665 0.610 ;
        RECT 1.215 0.270 1.385 0.415 ;
        RECT 2.105 0.085 2.475 0.580 ;
        RECT 3.325 0.085 3.595 0.720 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and2b_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__and2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and2b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 3.200 0.625 3.545 1.745 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.995 1.075 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.335 4.070 1.015 ;
        RECT 0.005 0.105 3.485 0.335 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.071500 ;
    PORT
      LAYER li1 ;
        RECT 1.635 1.535 2.980 1.745 ;
        RECT 2.445 0.825 2.980 1.535 ;
        RECT 1.675 0.615 2.980 0.825 ;
        RECT 1.675 0.495 1.865 0.615 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.090 2.255 0.425 2.635 ;
        RECT 1.090 2.275 1.420 2.635 ;
        RECT 2.055 2.275 2.435 2.635 ;
        RECT 2.995 2.275 3.375 2.635 ;
        RECT 0.165 1.915 3.940 2.085 ;
        RECT 0.165 1.325 0.335 1.915 ;
        RECT 0.515 1.500 1.415 1.745 ;
        RECT 1.245 1.485 1.415 1.500 ;
        RECT 1.245 1.355 1.420 1.485 ;
        RECT 0.165 0.995 0.425 1.325 ;
        RECT 1.245 0.995 2.175 1.355 ;
        RECT 1.245 0.805 1.455 0.995 ;
        RECT 0.090 0.615 1.455 0.805 ;
        RECT 0.090 0.255 0.425 0.615 ;
        RECT 3.725 0.495 3.940 1.915 ;
        RECT 1.055 0.085 1.385 0.445 ;
        RECT 2.035 0.085 2.415 0.445 ;
        RECT 2.995 0.085 3.375 0.445 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and2b_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__and3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.635 0.685 1.020 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.915 2.125 1.495 2.465 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.390 0.305 1.760 1.200 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.770 0.785 2.740 1.015 ;
        RECT 0.005 0.105 2.740 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 2.385 1.765 2.660 2.465 ;
        RECT 2.490 0.735 2.660 1.765 ;
        RECT 2.400 0.255 2.660 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.085 2.080 0.740 2.635 ;
        RECT 1.910 2.090 2.165 2.635 ;
        RECT 0.085 1.980 0.750 2.080 ;
        RECT 0.515 1.955 0.750 1.980 ;
        RECT 0.085 1.360 0.345 1.810 ;
        RECT 0.515 1.710 0.895 1.955 ;
        RECT 1.160 1.590 2.165 1.885 ;
        RECT 1.160 1.540 2.270 1.590 ;
        RECT 0.895 1.370 2.270 1.540 ;
        RECT 0.895 1.360 1.075 1.370 ;
        RECT 0.085 1.190 1.075 1.360 ;
        RECT 0.855 0.465 1.075 1.190 ;
        RECT 2.040 0.990 2.270 1.370 ;
        RECT 0.085 0.295 1.075 0.465 ;
        RECT 1.930 0.085 2.100 0.625 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and3_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__and3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.470 1.245 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.945 2.125 1.520 2.465 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.065 0.750 1.625 1.245 ;
        RECT 1.065 0.305 1.315 0.750 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.495 0.815 3.050 1.015 ;
        RECT 0.020 0.135 3.050 0.815 ;
        RECT 0.145 -0.085 0.315 0.135 ;
        RECT 1.510 0.105 3.050 0.135 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.511000 ;
    PORT
      LAYER li1 ;
        RECT 2.170 1.795 2.620 2.465 ;
        RECT 2.260 1.445 2.620 1.795 ;
        RECT 2.260 0.925 2.925 1.445 ;
        RECT 2.260 0.715 2.430 0.925 ;
        RECT 1.985 0.255 2.430 0.715 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.085 2.130 0.765 2.635 ;
        RECT 0.100 1.595 0.355 1.960 ;
        RECT 0.525 1.955 0.765 2.130 ;
        RECT 0.525 1.765 0.905 1.955 ;
        RECT 1.180 1.595 1.480 1.890 ;
        RECT 1.705 1.790 1.920 2.635 ;
        RECT 2.790 1.625 3.050 2.635 ;
        RECT 0.100 1.425 2.040 1.595 ;
        RECT 0.690 0.570 0.895 1.425 ;
        RECT 1.810 0.995 2.040 1.425 ;
        RECT 0.105 0.305 0.895 0.570 ;
        RECT 1.485 0.085 1.815 0.580 ;
        RECT 2.695 0.085 2.970 0.745 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and3_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__and3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.340 0.330 2.335 ;
        RECT 0.115 0.995 0.875 1.340 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.045 0.745 1.355 1.340 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.525 0.995 2.050 1.325 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.061500 ;
    PORT
      LAYER li1 ;
        RECT 2.650 1.760 2.840 2.465 ;
        RECT 3.610 1.765 3.800 2.465 ;
        RECT 3.610 1.760 4.490 1.765 ;
        RECT 2.650 1.535 4.490 1.760 ;
        RECT 4.210 0.845 4.490 1.535 ;
        RECT 2.650 0.615 4.490 0.845 ;
        RECT 2.650 0.515 2.840 0.615 ;
        RECT 3.610 0.255 3.800 0.615 ;
    END
  END X
  OBS
      LAYER pwell ;
        RECT 0.340 0.105 4.460 1.015 ;
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.500 1.750 0.680 2.465 ;
        RECT 0.895 1.935 1.395 2.635 ;
        RECT 1.620 1.750 1.800 2.465 ;
        RECT 2.060 1.935 2.390 2.635 ;
        RECT 3.010 1.935 3.390 2.635 ;
        RECT 3.970 1.935 4.350 2.635 ;
        RECT 0.500 1.580 2.430 1.750 ;
        RECT 2.220 1.355 2.430 1.580 ;
        RECT 2.220 1.020 3.905 1.355 ;
        RECT 2.220 0.805 2.430 1.020 ;
        RECT 0.465 0.445 0.800 0.805 ;
        RECT 1.635 0.615 2.430 0.805 ;
        RECT 1.635 0.445 1.825 0.615 ;
        RECT 0.465 0.255 1.825 0.445 ;
        RECT 2.055 0.085 2.385 0.445 ;
        RECT 3.010 0.085 3.390 0.445 ;
        RECT 3.970 0.085 4.350 0.445 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and3_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__and3b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and3b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.425 1.955 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.920 2.125 2.495 2.465 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 2.280 0.305 2.645 1.255 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.815 0.985 1.015 ;
        RECT 2.615 0.815 3.625 1.015 ;
        RECT 0.005 0.335 3.625 0.815 ;
        RECT 0.150 0.135 3.625 0.335 ;
        RECT 0.150 -0.085 0.320 0.135 ;
        RECT 2.630 0.105 3.625 0.135 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 3.270 1.765 3.535 2.465 ;
        RECT 3.365 0.735 3.535 1.765 ;
        RECT 3.275 0.255 3.535 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.085 2.125 0.345 2.635 ;
        RECT 0.645 1.245 0.815 2.465 ;
        RECT 1.085 2.130 1.750 2.635 ;
        RECT 1.505 1.955 1.750 2.130 ;
        RECT 2.795 2.090 3.010 2.635 ;
        RECT 1.085 1.595 1.335 1.940 ;
        RECT 1.505 1.765 1.885 1.955 ;
        RECT 2.155 1.595 3.050 1.890 ;
        RECT 1.085 1.575 3.050 1.595 ;
        RECT 1.085 1.425 3.185 1.575 ;
        RECT 0.645 0.995 1.520 1.245 ;
        RECT 0.645 0.905 0.895 0.995 ;
        RECT 0.085 0.085 0.345 0.905 ;
        RECT 0.515 0.485 0.895 0.905 ;
        RECT 1.690 0.550 1.945 1.425 ;
        RECT 2.965 0.975 3.185 1.425 ;
        RECT 1.105 0.285 1.945 0.550 ;
        RECT 2.815 0.085 3.105 0.625 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and3b_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__and3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and3b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.745 0.410 1.325 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.915 2.125 2.490 2.465 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.985 0.765 2.620 1.245 ;
        RECT 1.985 0.305 2.370 0.765 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.490 0.815 4.105 1.015 ;
        RECT 0.005 0.135 4.105 0.815 ;
        RECT 0.145 -0.085 0.315 0.135 ;
        RECT 2.505 0.105 4.105 0.135 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.498000 ;
    PORT
      LAYER li1 ;
        RECT 3.125 1.795 3.590 2.465 ;
        RECT 3.240 1.445 3.590 1.795 ;
        RECT 3.240 0.925 4.040 1.445 ;
        RECT 3.240 0.715 3.570 0.925 ;
        RECT 3.165 0.255 3.570 0.715 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.085 1.575 0.400 2.635 ;
        RECT 1.080 2.130 1.745 2.635 ;
        RECT 0.630 1.245 0.905 1.905 ;
        RECT 1.100 1.595 1.335 1.960 ;
        RECT 1.505 1.955 1.745 2.130 ;
        RECT 1.505 1.765 1.885 1.955 ;
        RECT 2.160 1.595 2.350 1.890 ;
        RECT 2.660 1.790 2.875 2.635 ;
        RECT 3.760 1.625 4.025 2.635 ;
        RECT 1.100 1.425 3.020 1.595 ;
        RECT 0.630 1.015 1.465 1.245 ;
        RECT 0.085 0.085 0.355 0.575 ;
        RECT 0.630 0.305 0.905 1.015 ;
        RECT 1.645 0.570 1.815 1.425 ;
        RECT 2.790 0.995 3.020 1.425 ;
        RECT 1.105 0.305 1.815 0.570 ;
        RECT 2.610 0.085 2.940 0.580 ;
        RECT 3.760 0.085 4.025 0.745 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and3b_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__and3b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and3b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 4.165 0.615 4.455 1.705 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.035 0.725 1.285 1.340 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.490 0.995 1.865 1.340 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.175 0.335 4.985 1.015 ;
        RECT 0.175 0.105 4.295 0.335 ;
        RECT 0.175 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.071500 ;
    PORT
      LAYER li1 ;
        RECT 2.375 1.535 3.995 1.705 ;
        RECT 3.570 0.845 3.995 1.535 ;
        RECT 2.485 0.615 3.995 0.845 ;
        RECT 2.485 0.515 2.675 0.615 ;
        RECT 3.365 0.255 3.635 0.615 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.060 2.805 ;
        RECT 0.730 2.275 1.230 2.635 ;
        RECT 1.895 2.275 2.225 2.635 ;
        RECT 2.845 2.275 3.230 2.635 ;
        RECT 3.805 2.275 4.185 2.635 ;
        RECT 0.150 1.495 0.510 2.165 ;
        RECT 0.680 1.875 4.905 2.105 ;
        RECT 0.150 0.805 0.370 1.495 ;
        RECT 0.680 1.325 0.865 1.875 ;
        RECT 1.330 1.525 2.205 1.695 ;
        RECT 0.540 0.995 0.865 1.325 ;
        RECT 2.035 1.355 2.205 1.525 ;
        RECT 2.035 1.020 3.400 1.355 ;
        RECT 2.035 0.805 2.265 1.020 ;
        RECT 0.150 0.545 0.635 0.805 ;
        RECT 1.520 0.615 2.265 0.805 ;
        RECT 1.520 0.545 1.700 0.615 ;
        RECT 0.150 0.355 1.700 0.545 ;
        RECT 0.150 0.255 0.635 0.355 ;
        RECT 1.930 0.085 2.260 0.445 ;
        RECT 2.845 0.085 3.195 0.445 ;
        RECT 3.805 0.085 4.185 0.445 ;
        RECT 4.625 0.425 4.905 1.875 ;
        RECT 0.000 -0.085 5.060 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and3b_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__and4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.325 2.075 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.855 0.360 1.235 1.325 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.405 0.355 1.695 1.325 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.885 0.715 2.165 1.325 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.930 0.785 3.165 1.015 ;
        RECT 0.005 0.105 3.165 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.752500 ;
    PORT
      LAYER li1 ;
        RECT 2.695 2.205 3.085 2.465 ;
        RECT 2.825 0.805 3.085 2.205 ;
        RECT 2.695 0.295 3.085 0.805 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.090 2.255 0.425 2.635 ;
        RECT 0.605 1.665 0.855 2.465 ;
        RECT 1.035 1.915 1.365 2.635 ;
        RECT 1.560 1.665 1.810 2.465 ;
        RECT 2.005 1.835 2.375 2.635 ;
        RECT 0.495 1.495 2.535 1.665 ;
        RECT 0.495 0.585 0.685 1.495 ;
        RECT 2.335 0.995 2.535 1.495 ;
        RECT 0.170 0.255 0.685 0.585 ;
        RECT 2.065 0.085 2.335 0.545 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and4_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__and4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.755 0.330 2.075 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.855 0.420 1.235 1.325 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.405 0.415 1.705 1.325 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.885 0.740 2.155 1.325 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.930 0.785 3.665 1.015 ;
        RECT 0.005 0.105 3.665 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.629500 ;
    PORT
      LAYER li1 ;
        RECT 2.625 1.835 3.075 2.465 ;
        RECT 2.835 0.805 3.075 1.835 ;
        RECT 2.625 0.295 3.075 0.805 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.095 2.255 0.425 2.635 ;
        RECT 0.645 1.665 0.815 2.465 ;
        RECT 1.035 1.915 1.365 2.635 ;
        RECT 1.570 1.665 1.820 2.465 ;
        RECT 2.165 1.835 2.415 2.635 ;
        RECT 3.245 1.835 3.565 2.635 ;
        RECT 0.500 1.495 2.665 1.665 ;
        RECT 0.500 0.585 0.670 1.495 ;
        RECT 2.495 0.995 2.665 1.495 ;
        RECT 0.175 0.255 0.670 0.585 ;
        RECT 2.285 0.085 2.455 0.550 ;
        RECT 3.245 0.085 3.575 0.810 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and4_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__and4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.765 0.330 1.655 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.890 0.420 1.345 1.325 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.515 0.425 1.780 1.325 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.985 0.730 2.275 1.325 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.535 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.028500 ;
    PORT
      LAYER li1 ;
        RECT 2.785 1.655 3.035 2.465 ;
        RECT 3.725 1.745 3.895 2.465 ;
        RECT 3.725 1.655 4.455 1.745 ;
        RECT 2.785 1.485 4.455 1.655 ;
        RECT 4.200 0.810 4.455 1.485 ;
        RECT 2.785 0.640 4.455 0.810 ;
        RECT 2.785 0.255 2.955 0.640 ;
        RECT 3.725 0.255 3.895 0.640 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.105 1.835 0.385 2.635 ;
        RECT 0.605 1.665 0.815 2.465 ;
        RECT 1.055 1.935 1.385 2.635 ;
        RECT 1.605 1.665 1.795 2.465 ;
        RECT 2.225 1.855 2.555 2.635 ;
        RECT 3.255 1.835 3.505 2.635 ;
        RECT 4.065 1.915 4.445 2.635 ;
        RECT 0.500 1.495 2.615 1.665 ;
        RECT 0.500 0.585 0.720 1.495 ;
        RECT 2.445 1.305 2.615 1.495 ;
        RECT 2.445 1.075 3.935 1.305 ;
        RECT 0.175 0.255 0.720 0.585 ;
        RECT 2.225 0.085 2.535 0.550 ;
        RECT 3.125 0.085 3.505 0.470 ;
        RECT 4.065 0.085 4.445 0.470 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and4_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__and4b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and4b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.450 1.675 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.675 0.420 2.155 1.695 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 2.325 0.420 2.615 1.695 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 2.785 0.665 3.075 1.695 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.995 0.785 3.975 1.015 ;
        RECT 0.005 0.105 3.975 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 3.635 1.495 3.995 2.465 ;
        RECT 3.725 0.805 3.995 1.495 ;
        RECT 3.520 0.295 3.995 0.805 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.170 2.015 0.345 2.465 ;
        RECT 0.515 2.195 0.895 2.635 ;
        RECT 1.200 2.045 1.370 2.465 ;
        RECT 1.655 2.225 2.375 2.635 ;
        RECT 2.630 2.045 2.800 2.465 ;
        RECT 3.060 2.225 3.390 2.635 ;
        RECT 0.170 1.845 0.850 2.015 ;
        RECT 0.680 1.325 0.850 1.845 ;
        RECT 1.200 1.875 3.415 2.045 ;
        RECT 0.680 0.995 1.025 1.325 ;
        RECT 0.680 0.825 0.850 0.995 ;
        RECT 0.170 0.655 0.850 0.825 ;
        RECT 0.170 0.255 0.345 0.655 ;
        RECT 1.200 0.585 1.370 1.875 ;
        RECT 3.245 1.325 3.415 1.875 ;
        RECT 3.245 0.995 3.535 1.325 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.140 0.255 1.370 0.585 ;
        RECT 2.955 0.085 3.350 0.465 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and4b_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__and4b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and4b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.135 0.740 0.335 1.630 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.895 0.420 2.155 1.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 2.375 0.420 2.615 1.615 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 2.785 0.645 3.115 1.615 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.045 0.785 4.535 1.015 ;
        RECT 0.005 0.105 4.535 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.555750 ;
    PORT
      LAYER li1 ;
        RECT 3.690 1.665 3.995 2.465 ;
        RECT 3.690 1.535 4.455 1.665 ;
        RECT 3.775 0.825 4.455 1.535 ;
        RECT 3.560 0.640 4.455 0.825 ;
        RECT 3.560 0.255 3.895 0.640 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.175 2.000 0.345 2.465 ;
        RECT 0.515 2.195 0.895 2.635 ;
        RECT 1.115 2.085 1.285 2.465 ;
        RECT 1.705 2.255 2.425 2.635 ;
        RECT 2.670 2.085 2.860 2.465 ;
        RECT 3.140 2.195 3.470 2.635 ;
        RECT 0.175 1.830 0.855 2.000 ;
        RECT 0.685 1.325 0.855 1.830 ;
        RECT 1.115 1.965 2.860 2.085 ;
        RECT 1.115 1.915 3.465 1.965 ;
        RECT 1.115 1.660 1.415 1.915 ;
        RECT 2.690 1.795 3.465 1.915 ;
        RECT 4.195 1.835 4.450 2.635 ;
        RECT 0.685 0.995 1.075 1.325 ;
        RECT 0.685 0.585 0.855 0.995 ;
        RECT 1.245 0.585 1.415 1.660 ;
        RECT 3.295 1.325 3.465 1.795 ;
        RECT 3.295 0.995 3.555 1.325 ;
        RECT 0.095 0.085 0.425 0.465 ;
        RECT 0.645 0.255 0.855 0.585 ;
        RECT 1.195 0.255 1.415 0.585 ;
        RECT 3.010 0.085 3.390 0.465 ;
        RECT 4.065 0.085 4.450 0.465 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and4b_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__and4b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and4b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.440 0.765 0.840 1.635 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 3.810 0.735 4.190 1.325 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 3.330 0.755 3.640 1.325 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.870 0.995 3.120 1.325 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.540 0.785 4.990 1.015 ;
        RECT 0.005 0.105 4.990 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.996000 ;
    PORT
      LAYER li1 ;
        RECT 1.030 1.545 2.360 1.715 ;
        RECT 1.030 0.820 1.360 1.545 ;
        RECT 1.030 0.650 2.280 0.820 ;
        RECT 1.030 0.255 1.340 0.650 ;
        RECT 2.110 0.255 2.280 0.650 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.060 2.805 ;
        RECT 0.085 2.085 0.345 2.465 ;
        RECT 0.515 2.255 0.895 2.635 ;
        RECT 1.510 2.255 1.890 2.635 ;
        RECT 2.450 2.255 2.830 2.635 ;
        RECT 3.510 2.255 3.890 2.635 ;
        RECT 4.570 2.255 4.950 2.635 ;
        RECT 0.085 1.915 4.885 2.085 ;
        RECT 0.085 0.585 0.260 1.915 ;
        RECT 2.530 1.545 4.530 1.715 ;
        RECT 2.530 1.325 2.700 1.545 ;
        RECT 1.530 0.995 2.700 1.325 ;
        RECT 4.360 0.810 4.530 1.545 ;
        RECT 4.715 0.995 4.885 1.915 ;
        RECT 4.360 0.640 4.900 0.810 ;
        RECT 0.085 0.255 0.345 0.585 ;
        RECT 0.565 0.085 0.815 0.545 ;
        RECT 1.510 0.085 1.890 0.470 ;
        RECT 2.535 0.085 2.865 0.445 ;
        RECT 0.000 -0.085 5.060 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and4b_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__and4bb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and4bb_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.625 0.815 1.955 ;
    END
  END A_N
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.525 0.945 1.165 1.115 ;
        RECT 0.525 0.765 0.785 0.945 ;
    END
  END B_N
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 2.875 0.415 3.175 1.635 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 3.345 0.420 3.640 1.635 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.565 0.785 4.590 1.015 ;
        RECT 0.005 0.335 4.590 0.785 ;
        RECT 0.005 0.105 1.525 0.335 ;
        RECT 3.620 0.105 4.590 0.335 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 4.250 1.445 4.510 2.465 ;
        RECT 4.285 0.825 4.510 1.445 ;
        RECT 4.250 0.255 4.510 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.085 2.135 0.345 2.465 ;
        RECT 0.575 2.255 0.955 2.635 ;
        RECT 0.085 1.455 0.255 2.135 ;
        RECT 1.165 2.085 1.375 2.465 ;
        RECT 1.625 2.255 1.955 2.635 ;
        RECT 2.185 2.085 2.355 2.465 ;
        RECT 2.550 2.255 2.930 2.635 ;
        RECT 3.210 2.085 3.380 2.465 ;
        RECT 3.700 2.255 4.030 2.635 ;
        RECT 1.165 1.915 1.985 2.085 ;
        RECT 1.015 1.575 1.645 1.745 ;
        RECT 1.015 1.455 1.235 1.575 ;
        RECT 0.085 1.285 1.235 1.455 ;
        RECT 1.815 1.405 1.985 1.915 ;
        RECT 0.085 0.585 0.255 1.285 ;
        RECT 1.415 1.235 1.985 1.405 ;
        RECT 2.155 1.915 3.980 2.085 ;
        RECT 1.415 0.755 1.585 1.235 ;
        RECT 2.155 0.925 2.325 1.915 ;
        RECT 3.810 1.325 3.980 1.915 ;
        RECT 0.085 0.255 0.345 0.585 ;
        RECT 0.575 0.085 0.955 0.465 ;
        RECT 1.185 0.425 1.585 0.755 ;
        RECT 1.755 0.595 2.325 0.925 ;
        RECT 2.495 0.425 2.665 1.325 ;
        RECT 3.810 0.995 4.115 1.325 ;
        RECT 1.185 0.255 2.665 0.425 ;
        RECT 3.810 0.085 3.980 0.545 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and4bb_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__and4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and4bb_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.150 0.995 0.330 1.635 ;
    END
  END A_N
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 4.175 0.765 4.525 1.305 ;
    END
  END B_N
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 3.270 0.420 3.535 1.275 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 3.705 0.425 4.005 1.405 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.540 0.785 1.965 1.015 ;
        RECT 0.005 0.105 4.995 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.498000 ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.545 1.420 1.715 ;
        RECT 1.065 0.255 1.340 1.545 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.060 2.805 ;
        RECT 0.175 2.055 0.345 2.465 ;
        RECT 0.515 2.255 0.895 2.635 ;
        RECT 1.640 2.255 2.310 2.635 ;
        RECT 2.595 2.085 2.765 2.465 ;
        RECT 2.935 2.255 3.325 2.635 ;
        RECT 3.545 2.085 3.715 2.465 ;
        RECT 4.105 2.255 4.435 2.635 ;
        RECT 4.655 2.085 4.915 2.465 ;
        RECT 0.175 1.885 2.075 2.055 ;
        RECT 0.500 0.805 0.720 1.885 ;
        RECT 1.905 1.325 2.075 1.885 ;
        RECT 2.385 1.915 3.715 2.085 ;
        RECT 3.885 1.915 4.915 2.085 ;
        RECT 0.175 0.635 0.720 0.805 ;
        RECT 1.515 0.805 1.735 1.325 ;
        RECT 1.905 0.995 2.215 1.325 ;
        RECT 2.385 0.805 2.605 1.915 ;
        RECT 3.885 1.745 4.105 1.915 ;
        RECT 2.795 1.575 4.105 1.745 ;
        RECT 2.795 1.400 3.015 1.575 ;
        RECT 1.515 0.635 2.605 0.805 ;
        RECT 0.175 0.255 0.345 0.635 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.510 0.085 1.890 0.465 ;
        RECT 2.145 0.255 2.315 0.635 ;
        RECT 4.745 0.585 4.915 1.915 ;
        RECT 4.185 0.085 4.435 0.585 ;
        RECT 4.655 0.255 4.915 0.585 ;
        RECT 0.000 -0.085 5.060 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and4bb_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__and4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and4bb_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 5.935 0.995 6.345 1.620 ;
    END
  END A_N
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.430 0.765 0.830 1.635 ;
    END
  END B_N
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 3.365 0.640 3.840 1.325 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.905 0.995 3.195 1.325 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.540 0.785 5.150 1.015 ;
        RECT 0.005 0.105 6.435 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.996000 ;
    PORT
      LAYER li1 ;
        RECT 1.010 1.545 2.360 1.715 ;
        RECT 1.010 0.820 1.340 1.545 ;
        RECT 1.010 0.650 2.280 0.820 ;
        RECT 1.170 0.255 1.340 0.650 ;
        RECT 2.110 0.255 2.280 0.650 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.085 2.085 0.345 2.465 ;
        RECT 0.515 2.255 0.895 2.635 ;
        RECT 1.510 2.255 1.890 2.635 ;
        RECT 2.450 2.255 2.830 2.635 ;
        RECT 3.680 2.255 4.010 2.635 ;
        RECT 4.810 2.255 5.820 2.635 ;
        RECT 6.095 2.085 6.265 2.465 ;
        RECT 0.085 1.915 4.940 2.085 ;
        RECT 0.085 0.585 0.260 1.915 ;
        RECT 2.530 1.545 4.550 1.715 ;
        RECT 2.530 1.245 2.700 1.545 ;
        RECT 4.770 1.375 4.940 1.915 ;
        RECT 1.510 1.075 2.700 1.245 ;
        RECT 2.530 0.785 2.700 1.075 ;
        RECT 4.080 1.205 4.940 1.375 ;
        RECT 5.360 1.915 6.265 2.085 ;
        RECT 4.080 0.995 4.300 1.205 ;
        RECT 5.360 0.825 5.530 1.915 ;
        RECT 2.530 0.615 3.195 0.785 ;
        RECT 0.085 0.255 0.345 0.585 ;
        RECT 2.975 0.470 3.195 0.615 ;
        RECT 4.710 0.470 5.060 0.810 ;
        RECT 5.360 0.655 6.265 0.825 ;
        RECT 0.620 0.085 0.950 0.470 ;
        RECT 1.510 0.085 1.890 0.470 ;
        RECT 2.470 0.085 2.800 0.445 ;
        RECT 2.975 0.300 5.060 0.470 ;
        RECT 5.385 0.085 5.715 0.465 ;
        RECT 6.095 0.255 6.265 0.655 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and4bb_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__buf_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__buf_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.220200 ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.985 0.545 1.355 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 1.475 0.885 ;
        RECT 0.155 -0.085 0.325 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.348500 ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.560 1.395 2.465 ;
        RECT 1.215 0.760 1.395 1.560 ;
        RECT 1.065 0.255 1.395 0.760 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.840 2.805 ;
        RECT 0.165 1.705 0.345 2.465 ;
        RECT 0.525 1.875 0.895 2.635 ;
        RECT 0.165 1.535 0.890 1.705 ;
        RECT 0.720 1.390 0.890 1.535 ;
        RECT 0.720 1.060 1.035 1.390 ;
        RECT 0.720 0.805 0.890 1.060 ;
        RECT 0.175 0.635 0.890 0.805 ;
        RECT 0.175 0.255 0.345 0.635 ;
        RECT 0.525 0.085 0.895 0.465 ;
        RECT 0.000 -0.085 1.840 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__buf_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__buf_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__buf_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.440 1.355 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.540 0.785 2.210 1.015 ;
        RECT 0.005 0.105 2.210 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.703750 ;
    PORT
      LAYER li1 ;
        RECT 1.270 0.255 1.695 2.465 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.175 1.705 0.345 2.465 ;
        RECT 0.600 1.875 0.930 2.635 ;
        RECT 0.175 1.535 0.895 1.705 ;
        RECT 0.725 1.325 0.895 1.535 ;
        RECT 1.865 1.485 2.125 2.635 ;
        RECT 0.725 0.995 1.025 1.325 ;
        RECT 0.725 0.805 0.940 0.995 ;
        RECT 0.175 0.635 0.940 0.805 ;
        RECT 0.175 0.255 0.345 0.635 ;
        RECT 0.610 0.085 0.940 0.465 ;
        RECT 1.865 0.085 2.125 0.925 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__buf_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__buf_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__buf_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 0.470 1.315 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.865 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.996000 ;
    PORT
      LAYER li1 ;
        RECT 1.115 1.615 1.285 2.465 ;
        RECT 2.055 1.615 2.225 2.465 ;
        RECT 1.115 1.445 2.225 1.615 ;
        RECT 1.920 0.905 2.225 1.445 ;
        RECT 1.115 0.735 2.225 0.905 ;
        RECT 1.115 0.255 1.285 0.735 ;
        RECT 2.055 0.255 2.225 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.095 1.655 0.425 2.465 ;
        RECT 0.645 1.835 0.885 2.635 ;
        RECT 1.455 1.835 1.835 2.635 ;
        RECT 0.095 1.485 0.860 1.655 ;
        RECT 2.395 1.485 2.775 2.635 ;
        RECT 0.690 1.245 0.860 1.485 ;
        RECT 0.690 1.075 1.240 1.245 ;
        RECT 0.690 0.905 0.860 1.075 ;
        RECT 0.175 0.735 0.860 0.905 ;
        RECT 0.175 0.255 0.345 0.735 ;
        RECT 0.525 0.085 0.815 0.565 ;
        RECT 1.455 0.085 1.835 0.565 ;
        RECT 2.395 0.085 2.775 0.885 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__buf_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__buf_6
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__buf_6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.280 1.075 1.265 1.315 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.265 0.105 4.535 1.015 ;
        RECT 0.265 0.085 0.320 0.105 ;
        RECT 0.150 -0.085 0.320 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.526500 ;
    PORT
      LAYER li1 ;
        RECT 1.845 1.615 2.015 2.465 ;
        RECT 2.785 1.615 2.955 2.465 ;
        RECT 3.725 1.615 3.895 2.465 ;
        RECT 1.845 1.445 3.895 1.615 ;
        RECT 2.410 0.905 3.895 1.445 ;
        RECT 1.845 0.735 3.895 0.905 ;
        RECT 1.845 0.255 2.015 0.735 ;
        RECT 2.785 0.255 2.955 0.735 ;
        RECT 3.725 0.255 3.895 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.435 1.485 0.605 2.635 ;
        RECT 0.775 1.655 1.155 2.465 ;
        RECT 1.375 1.835 1.615 2.635 ;
        RECT 2.185 1.835 2.565 2.635 ;
        RECT 3.125 1.835 3.505 2.635 ;
        RECT 0.775 1.485 1.625 1.655 ;
        RECT 4.065 1.485 4.445 2.635 ;
        RECT 1.455 1.245 1.625 1.485 ;
        RECT 1.455 1.075 1.975 1.245 ;
        RECT 1.455 0.905 1.625 1.075 ;
        RECT 0.775 0.735 1.625 0.905 ;
        RECT 0.435 0.085 0.605 0.565 ;
        RECT 0.775 0.255 1.155 0.735 ;
        RECT 1.375 0.085 1.545 0.565 ;
        RECT 2.185 0.085 2.565 0.565 ;
        RECT 3.125 0.085 3.505 0.565 ;
        RECT 4.065 0.085 4.445 0.885 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__buf_6

#--------EOF---------

MACRO sky130_fd_sc_hdll__buf_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__buf_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.832500 ;
    PORT
      LAYER li1 ;
        RECT 0.140 1.075 1.340 1.275 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.685 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.024500 ;
    PORT
      LAYER li1 ;
        RECT 2.055 1.615 2.225 2.465 ;
        RECT 2.995 1.615 3.165 2.465 ;
        RECT 3.935 1.615 4.105 2.465 ;
        RECT 4.875 1.615 5.045 2.465 ;
        RECT 2.055 1.445 5.045 1.615 ;
        RECT 4.690 0.905 5.045 1.445 ;
        RECT 2.055 0.735 5.045 0.905 ;
        RECT 2.055 0.255 2.225 0.735 ;
        RECT 2.995 0.255 3.165 0.735 ;
        RECT 3.935 0.255 4.105 0.735 ;
        RECT 4.875 0.255 5.045 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.095 1.615 0.425 2.465 ;
        RECT 0.645 1.835 0.815 2.635 ;
        RECT 0.985 1.615 1.365 2.465 ;
        RECT 1.585 1.835 1.755 2.635 ;
        RECT 2.395 1.835 2.775 2.635 ;
        RECT 3.335 1.835 3.715 2.635 ;
        RECT 4.275 1.835 4.655 2.635 ;
        RECT 0.095 1.445 1.745 1.615 ;
        RECT 5.215 1.485 5.595 2.635 ;
        RECT 1.570 1.245 1.745 1.445 ;
        RECT 1.570 1.075 4.495 1.245 ;
        RECT 1.570 0.905 1.745 1.075 ;
        RECT 0.175 0.735 1.745 0.905 ;
        RECT 0.175 0.255 0.345 0.735 ;
        RECT 0.515 0.085 0.895 0.565 ;
        RECT 1.115 0.260 1.285 0.735 ;
        RECT 1.455 0.085 1.835 0.565 ;
        RECT 2.395 0.085 2.775 0.565 ;
        RECT 3.335 0.085 3.715 0.565 ;
        RECT 4.275 0.085 4.655 0.565 ;
        RECT 5.215 0.085 5.595 0.885 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__buf_8

#--------EOF---------

MACRO sky130_fd_sc_hdll__buf_12
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__buf_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.280 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.135 1.075 1.810 1.275 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.280 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 8.075 1.015 ;
        RECT 0.620 -0.085 0.790 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.470 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.280 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.020500 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.615 2.695 2.465 ;
        RECT 3.465 1.615 3.635 2.465 ;
        RECT 4.405 1.615 4.575 2.465 ;
        RECT 5.345 1.615 5.515 2.465 ;
        RECT 6.285 1.615 6.455 2.465 ;
        RECT 7.225 1.615 7.395 2.465 ;
        RECT 2.525 1.445 7.395 1.615 ;
        RECT 5.210 0.905 7.395 1.445 ;
        RECT 2.525 0.735 7.395 0.905 ;
        RECT 2.525 0.255 2.695 0.735 ;
        RECT 3.465 0.255 3.635 0.735 ;
        RECT 4.405 0.255 4.575 0.735 ;
        RECT 5.345 0.255 5.515 0.735 ;
        RECT 6.285 0.255 6.455 0.735 ;
        RECT 7.225 0.255 7.395 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.280 2.805 ;
        RECT 0.175 1.835 0.345 2.635 ;
        RECT 0.515 1.615 0.895 2.465 ;
        RECT 1.115 1.835 1.285 2.635 ;
        RECT 1.455 1.615 1.835 2.465 ;
        RECT 2.055 1.835 2.225 2.635 ;
        RECT 2.865 1.835 3.245 2.635 ;
        RECT 3.805 1.835 4.185 2.635 ;
        RECT 4.745 1.835 5.125 2.635 ;
        RECT 5.685 1.835 6.065 2.635 ;
        RECT 6.625 1.835 7.005 2.635 ;
        RECT 0.515 1.445 2.215 1.615 ;
        RECT 7.565 1.485 7.945 2.635 ;
        RECT 2.040 1.245 2.215 1.445 ;
        RECT 2.040 1.075 4.965 1.245 ;
        RECT 2.040 0.905 2.215 1.075 ;
        RECT 0.645 0.735 2.215 0.905 ;
        RECT 0.095 0.085 0.425 0.565 ;
        RECT 0.645 0.255 0.815 0.735 ;
        RECT 0.985 0.085 1.365 0.565 ;
        RECT 1.585 0.260 1.755 0.735 ;
        RECT 1.925 0.085 2.305 0.565 ;
        RECT 2.865 0.085 3.245 0.565 ;
        RECT 3.805 0.085 4.185 0.565 ;
        RECT 4.745 0.085 5.125 0.565 ;
        RECT 5.685 0.085 6.065 0.565 ;
        RECT 6.625 0.085 7.005 0.565 ;
        RECT 7.565 0.085 7.945 0.885 ;
        RECT 0.000 -0.085 8.280 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__buf_12

#--------EOF---------

MACRO sky130_fd_sc_hdll__buf_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__buf_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.500 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.665000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 2.735 1.275 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.500 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 10.855 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 11.690 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.500 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.016500 ;
    PORT
      LAYER li1 ;
        RECT 3.335 1.615 3.715 2.465 ;
        RECT 4.275 1.615 4.655 2.465 ;
        RECT 5.215 1.615 5.595 2.465 ;
        RECT 6.155 1.615 6.535 2.465 ;
        RECT 7.095 1.615 7.475 2.465 ;
        RECT 8.035 1.615 8.415 2.465 ;
        RECT 8.975 1.615 9.355 2.465 ;
        RECT 9.915 1.615 10.295 2.465 ;
        RECT 10.860 1.615 11.135 2.360 ;
        RECT 3.335 1.445 11.135 1.615 ;
        RECT 10.635 0.905 11.135 1.445 ;
        RECT 3.335 0.735 11.135 0.905 ;
        RECT 3.335 0.260 3.715 0.735 ;
        RECT 4.275 0.260 4.655 0.735 ;
        RECT 5.215 0.260 5.595 0.735 ;
        RECT 6.155 0.260 6.535 0.735 ;
        RECT 7.095 0.260 7.475 0.735 ;
        RECT 8.035 0.260 8.415 0.735 ;
        RECT 8.975 0.260 9.355 0.735 ;
        RECT 9.915 0.260 10.295 0.735 ;
        RECT 10.860 0.365 11.135 0.735 ;
        RECT 3.335 0.255 3.635 0.260 ;
        RECT 4.405 0.255 4.575 0.260 ;
        RECT 5.345 0.255 5.515 0.260 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 11.500 2.805 ;
        RECT 0.175 1.445 0.345 2.635 ;
        RECT 0.515 1.615 0.895 2.465 ;
        RECT 1.115 1.835 1.285 2.635 ;
        RECT 1.455 1.615 1.835 2.465 ;
        RECT 2.055 1.835 2.225 2.635 ;
        RECT 2.395 1.615 2.775 2.465 ;
        RECT 2.995 1.835 3.165 2.635 ;
        RECT 3.935 1.835 4.105 2.635 ;
        RECT 4.875 1.835 5.045 2.635 ;
        RECT 5.815 1.835 5.985 2.635 ;
        RECT 6.755 1.835 6.925 2.635 ;
        RECT 7.695 1.835 7.865 2.635 ;
        RECT 8.635 1.835 8.805 2.635 ;
        RECT 9.575 1.835 9.745 2.635 ;
        RECT 10.515 1.835 10.685 2.635 ;
        RECT 0.515 1.445 3.165 1.615 ;
        RECT 2.990 1.275 3.165 1.445 ;
        RECT 2.990 1.075 10.175 1.275 ;
        RECT 2.990 0.905 3.165 1.075 ;
        RECT 0.175 0.085 0.345 0.905 ;
        RECT 0.515 0.735 3.165 0.905 ;
        RECT 0.515 0.260 0.895 0.735 ;
        RECT 1.115 0.085 1.285 0.565 ;
        RECT 1.455 0.260 1.835 0.735 ;
        RECT 2.055 0.085 2.225 0.565 ;
        RECT 2.395 0.260 2.775 0.735 ;
        RECT 2.995 0.085 3.165 0.565 ;
        RECT 3.935 0.085 4.105 0.565 ;
        RECT 4.875 0.085 5.045 0.565 ;
        RECT 5.815 0.085 5.985 0.565 ;
        RECT 6.755 0.085 6.925 0.565 ;
        RECT 7.695 0.085 7.865 0.565 ;
        RECT 8.635 0.085 8.805 0.565 ;
        RECT 9.575 0.085 9.745 0.565 ;
        RECT 10.515 0.085 10.685 0.565 ;
        RECT 0.000 -0.085 11.500 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__buf_16

#--------EOF---------

MACRO sky130_fd_sc_hdll__bufbuf_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__bufbuf_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.110 1.075 0.440 1.275 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.540 0.785 7.240 1.015 ;
        RECT 0.005 0.105 7.240 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.024500 ;
    PORT
      LAYER li1 ;
        RECT 3.480 1.615 3.860 2.465 ;
        RECT 4.420 1.615 4.800 2.465 ;
        RECT 5.360 1.615 5.740 2.465 ;
        RECT 6.300 1.615 6.680 2.465 ;
        RECT 3.480 1.445 7.240 1.615 ;
        RECT 6.860 0.905 7.240 1.445 ;
        RECT 3.480 0.735 7.240 0.905 ;
        RECT 3.480 0.260 3.860 0.735 ;
        RECT 4.420 0.260 4.800 0.735 ;
        RECT 5.360 0.260 5.740 0.735 ;
        RECT 6.300 0.260 6.680 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.360 2.805 ;
        RECT 0.095 1.615 0.425 2.160 ;
        RECT 0.645 1.785 0.815 2.635 ;
        RECT 0.095 1.445 0.830 1.615 ;
        RECT 1.050 1.545 1.480 2.465 ;
        RECT 0.660 1.325 0.830 1.445 ;
        RECT 0.660 0.995 1.140 1.325 ;
        RECT 1.310 1.275 1.480 1.545 ;
        RECT 1.650 1.615 1.980 2.465 ;
        RECT 2.200 1.785 2.370 2.635 ;
        RECT 2.540 1.615 2.920 2.465 ;
        RECT 3.140 1.785 3.310 2.635 ;
        RECT 4.080 1.835 4.250 2.635 ;
        RECT 5.020 1.835 5.190 2.635 ;
        RECT 5.960 1.835 6.130 2.635 ;
        RECT 6.900 1.835 7.070 2.635 ;
        RECT 1.650 1.445 3.310 1.615 ;
        RECT 3.140 1.275 3.310 1.445 ;
        RECT 1.310 1.075 2.920 1.275 ;
        RECT 3.140 1.075 5.910 1.275 ;
        RECT 0.660 0.905 0.830 0.995 ;
        RECT 0.095 0.735 0.830 0.905 ;
        RECT 1.310 0.825 1.480 1.075 ;
        RECT 3.140 0.905 3.310 1.075 ;
        RECT 0.095 0.260 0.425 0.735 ;
        RECT 0.645 0.085 0.815 0.565 ;
        RECT 1.050 0.260 1.480 0.825 ;
        RECT 1.650 0.735 3.310 0.905 ;
        RECT 1.650 0.260 1.980 0.735 ;
        RECT 2.200 0.085 2.370 0.565 ;
        RECT 2.540 0.260 2.920 0.735 ;
        RECT 3.140 0.085 3.310 0.565 ;
        RECT 4.080 0.085 4.250 0.565 ;
        RECT 5.020 0.085 5.190 0.565 ;
        RECT 5.960 0.085 6.130 0.565 ;
        RECT 6.900 0.085 7.070 0.565 ;
        RECT 0.000 -0.085 7.360 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__bufbuf_8

#--------EOF---------

MACRO sky130_fd_sc_hdll__bufbuf_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__bufbuf_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.340 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.110 1.075 0.440 1.275 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 13.340 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 13.255 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 13.530 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 13.340 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.016500 ;
    PORT
      LAYER li1 ;
        RECT 5.735 1.615 6.115 2.465 ;
        RECT 6.675 1.615 7.055 2.465 ;
        RECT 7.615 1.615 7.995 2.465 ;
        RECT 8.555 1.615 8.935 2.465 ;
        RECT 9.495 1.615 9.875 2.465 ;
        RECT 10.435 1.615 10.815 2.465 ;
        RECT 11.375 1.615 11.755 2.465 ;
        RECT 12.315 1.615 12.695 2.465 ;
        RECT 5.735 1.445 13.220 1.615 ;
        RECT 12.920 0.905 13.220 1.445 ;
        RECT 5.735 0.735 13.220 0.905 ;
        RECT 5.735 0.260 6.115 0.735 ;
        RECT 6.675 0.260 7.055 0.735 ;
        RECT 7.615 0.260 7.995 0.735 ;
        RECT 8.555 0.260 8.935 0.735 ;
        RECT 9.495 0.260 9.875 0.735 ;
        RECT 10.435 0.260 10.815 0.735 ;
        RECT 11.375 0.260 11.755 0.735 ;
        RECT 12.315 0.260 12.695 0.735 ;
        RECT 5.735 0.255 6.035 0.260 ;
        RECT 6.805 0.255 6.975 0.260 ;
        RECT 7.745 0.255 7.915 0.260 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 13.340 2.805 ;
        RECT 0.175 1.445 0.345 2.635 ;
        RECT 0.515 1.445 0.895 2.465 ;
        RECT 1.085 1.615 1.415 2.465 ;
        RECT 1.635 1.785 1.805 2.635 ;
        RECT 1.975 1.615 2.355 2.465 ;
        RECT 2.575 1.785 2.745 2.635 ;
        RECT 2.915 1.615 3.295 2.465 ;
        RECT 3.515 1.835 3.685 2.635 ;
        RECT 3.855 1.615 4.235 2.465 ;
        RECT 4.455 1.835 4.625 2.635 ;
        RECT 4.795 1.615 5.175 2.465 ;
        RECT 5.395 1.835 5.565 2.635 ;
        RECT 6.335 1.835 6.505 2.635 ;
        RECT 7.275 1.835 7.445 2.635 ;
        RECT 8.215 1.835 8.385 2.635 ;
        RECT 9.155 1.835 9.325 2.635 ;
        RECT 10.095 1.835 10.265 2.635 ;
        RECT 11.035 1.835 11.205 2.635 ;
        RECT 11.975 1.835 12.145 2.635 ;
        RECT 12.915 1.835 13.085 2.635 ;
        RECT 1.085 1.445 2.745 1.615 ;
        RECT 2.915 1.445 5.565 1.615 ;
        RECT 0.660 1.275 0.895 1.445 ;
        RECT 2.575 1.275 2.745 1.445 ;
        RECT 5.390 1.275 5.565 1.445 ;
        RECT 0.660 1.075 2.355 1.275 ;
        RECT 2.575 1.075 5.135 1.275 ;
        RECT 5.390 1.075 12.700 1.275 ;
        RECT 0.660 0.905 0.895 1.075 ;
        RECT 2.575 0.905 2.745 1.075 ;
        RECT 5.390 0.905 5.565 1.075 ;
        RECT 0.175 0.085 0.345 0.905 ;
        RECT 0.515 0.260 0.895 0.905 ;
        RECT 1.085 0.735 2.745 0.905 ;
        RECT 2.915 0.735 5.565 0.905 ;
        RECT 1.085 0.260 1.415 0.735 ;
        RECT 1.635 0.085 1.805 0.565 ;
        RECT 1.975 0.260 2.355 0.735 ;
        RECT 2.575 0.085 2.745 0.565 ;
        RECT 2.915 0.260 3.295 0.735 ;
        RECT 3.515 0.085 3.685 0.565 ;
        RECT 3.855 0.260 4.235 0.735 ;
        RECT 4.455 0.085 4.625 0.565 ;
        RECT 4.795 0.260 5.175 0.735 ;
        RECT 5.395 0.085 5.565 0.565 ;
        RECT 6.335 0.085 6.505 0.565 ;
        RECT 7.275 0.085 7.445 0.565 ;
        RECT 8.215 0.085 8.385 0.565 ;
        RECT 9.155 0.085 9.325 0.565 ;
        RECT 10.095 0.085 10.265 0.565 ;
        RECT 11.035 0.085 11.205 0.565 ;
        RECT 11.975 0.085 12.145 0.565 ;
        RECT 12.915 0.085 13.085 0.565 ;
        RECT 0.000 -0.085 13.340 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__bufbuf_16

#--------EOF---------

MACRO sky130_fd_sc_hdll__bufinv_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__bufinv_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.900 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.505 1.275 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.900 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 6.675 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.090 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.900 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.024500 ;
    PORT
      LAYER li1 ;
        RECT 2.915 1.615 3.295 2.465 ;
        RECT 3.855 1.615 4.235 2.465 ;
        RECT 4.795 1.615 5.175 2.465 ;
        RECT 5.735 1.615 6.115 2.465 ;
        RECT 2.915 1.445 6.805 1.615 ;
        RECT 6.415 0.905 6.805 1.445 ;
        RECT 2.915 0.735 6.805 0.905 ;
        RECT 2.915 0.260 3.295 0.735 ;
        RECT 3.855 0.260 4.235 0.735 ;
        RECT 4.795 0.260 5.175 0.735 ;
        RECT 5.735 0.260 6.115 0.735 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.900 2.805 ;
        RECT 0.175 1.445 0.345 2.635 ;
        RECT 0.515 1.545 0.895 2.465 ;
        RECT 0.725 1.275 0.895 1.545 ;
        RECT 1.085 1.615 1.415 2.465 ;
        RECT 1.635 1.785 1.805 2.635 ;
        RECT 1.975 1.615 2.355 2.465 ;
        RECT 2.575 1.785 2.745 2.635 ;
        RECT 3.515 1.835 3.685 2.635 ;
        RECT 4.455 1.835 4.625 2.635 ;
        RECT 5.395 1.835 5.565 2.635 ;
        RECT 6.335 1.835 6.505 2.635 ;
        RECT 1.085 1.445 2.745 1.615 ;
        RECT 2.575 1.275 2.745 1.445 ;
        RECT 0.725 1.075 2.355 1.275 ;
        RECT 2.575 1.075 6.245 1.275 ;
        RECT 0.725 0.905 0.895 1.075 ;
        RECT 2.575 0.905 2.745 1.075 ;
        RECT 0.175 0.085 0.345 0.905 ;
        RECT 0.515 0.260 0.895 0.905 ;
        RECT 1.085 0.735 2.745 0.905 ;
        RECT 1.085 0.260 1.415 0.735 ;
        RECT 1.635 0.085 1.805 0.565 ;
        RECT 1.975 0.260 2.355 0.735 ;
        RECT 2.575 0.085 2.745 0.565 ;
        RECT 3.515 0.085 3.685 0.565 ;
        RECT 4.455 0.085 4.625 0.565 ;
        RECT 5.395 0.085 5.565 0.565 ;
        RECT 6.335 0.085 6.505 0.565 ;
        RECT 0.000 -0.085 6.900 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__bufinv_8

#--------EOF---------

MACRO sky130_fd_sc_hdll__bufinv_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__bufinv_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.420 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.832500 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 1.365 1.275 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 12.420 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 12.265 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 12.610 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 12.420 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.016500 ;
    PORT
      LAYER li1 ;
        RECT 4.745 1.615 5.125 2.465 ;
        RECT 5.685 1.615 6.065 2.465 ;
        RECT 6.625 1.615 7.005 2.465 ;
        RECT 7.565 1.615 7.945 2.465 ;
        RECT 8.505 1.615 8.885 2.465 ;
        RECT 9.445 1.615 9.825 2.465 ;
        RECT 10.385 1.615 10.765 2.465 ;
        RECT 11.325 1.615 11.705 2.465 ;
        RECT 4.745 1.445 12.205 1.615 ;
        RECT 11.930 0.905 12.205 1.445 ;
        RECT 4.745 0.735 12.205 0.905 ;
        RECT 4.745 0.260 5.125 0.735 ;
        RECT 5.685 0.260 6.065 0.735 ;
        RECT 6.625 0.260 7.005 0.735 ;
        RECT 7.565 0.260 7.945 0.735 ;
        RECT 8.505 0.260 8.885 0.735 ;
        RECT 9.445 0.260 9.825 0.735 ;
        RECT 10.385 0.260 10.765 0.735 ;
        RECT 11.325 0.260 11.705 0.735 ;
        RECT 4.745 0.255 5.045 0.260 ;
        RECT 5.815 0.255 5.985 0.260 ;
        RECT 6.755 0.255 6.925 0.260 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 12.420 2.805 ;
        RECT 0.095 1.615 0.425 2.465 ;
        RECT 0.645 1.785 0.815 2.635 ;
        RECT 0.985 1.615 1.365 2.465 ;
        RECT 1.585 1.785 1.755 2.635 ;
        RECT 1.925 1.615 2.305 2.465 ;
        RECT 2.525 1.835 2.695 2.635 ;
        RECT 2.865 1.615 3.245 2.465 ;
        RECT 3.465 1.835 3.635 2.635 ;
        RECT 3.805 1.615 4.185 2.465 ;
        RECT 4.405 1.835 4.575 2.635 ;
        RECT 5.345 1.835 5.515 2.635 ;
        RECT 6.285 1.835 6.455 2.635 ;
        RECT 7.225 1.835 7.395 2.635 ;
        RECT 8.165 1.835 8.335 2.635 ;
        RECT 9.105 1.835 9.275 2.635 ;
        RECT 10.045 1.835 10.215 2.635 ;
        RECT 10.985 1.835 11.155 2.635 ;
        RECT 11.925 1.835 12.095 2.635 ;
        RECT 0.095 1.445 1.755 1.615 ;
        RECT 1.925 1.445 4.575 1.615 ;
        RECT 1.585 1.275 1.755 1.445 ;
        RECT 4.400 1.275 4.575 1.445 ;
        RECT 1.585 1.075 4.145 1.275 ;
        RECT 4.400 1.075 11.710 1.275 ;
        RECT 1.585 0.905 1.755 1.075 ;
        RECT 4.400 0.905 4.575 1.075 ;
        RECT 0.095 0.735 1.755 0.905 ;
        RECT 1.925 0.735 4.575 0.905 ;
        RECT 0.095 0.260 0.425 0.735 ;
        RECT 0.645 0.085 0.815 0.565 ;
        RECT 0.985 0.260 1.365 0.735 ;
        RECT 1.585 0.085 1.755 0.565 ;
        RECT 1.925 0.260 2.305 0.735 ;
        RECT 2.525 0.085 2.695 0.565 ;
        RECT 2.865 0.260 3.245 0.735 ;
        RECT 3.465 0.085 3.635 0.565 ;
        RECT 3.805 0.260 4.185 0.735 ;
        RECT 4.405 0.085 4.575 0.565 ;
        RECT 5.345 0.085 5.515 0.565 ;
        RECT 6.285 0.085 6.455 0.565 ;
        RECT 7.225 0.085 7.395 0.565 ;
        RECT 8.165 0.085 8.335 0.565 ;
        RECT 9.105 0.085 9.275 0.565 ;
        RECT 10.045 0.085 10.215 0.565 ;
        RECT 10.985 0.085 11.155 0.565 ;
        RECT 11.925 0.085 12.095 0.565 ;
        RECT 0.000 -0.085 12.420 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__bufinv_16

#--------EOF---------

MACRO sky130_fd_sc_hdll__clkbuf_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__clkbuf_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.220200 ;
    PORT
      LAYER li1 ;
        RECT 1.365 0.985 1.745 1.355 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VPB
    DIRECTION INPUT ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.374500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.560 0.355 2.465 ;
        RECT 0.085 0.760 0.255 1.560 ;
        RECT 0.085 0.255 0.345 0.760 ;
    END
  END X
  OBS
      LAYER pwell ;
        RECT 0.005 0.105 1.795 0.885 ;
        RECT 1.165 -0.085 1.335 0.105 ;
      LAYER li1 ;
        RECT 0.000 2.635 1.840 2.805 ;
        RECT 0.525 1.875 1.275 2.635 ;
        RECT 1.495 1.705 1.665 2.465 ;
        RECT 0.540 1.535 1.665 1.705 ;
        RECT 0.540 1.390 0.760 1.535 ;
        RECT 0.425 1.060 0.760 1.390 ;
        RECT 0.540 0.805 0.760 1.060 ;
        RECT 0.540 0.635 1.625 0.805 ;
        RECT 0.525 0.085 1.275 0.465 ;
        RECT 1.455 0.255 1.625 0.635 ;
        RECT 0.000 -0.085 1.840 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkbuf_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__clkbuf_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__clkbuf_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.243000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.745 0.835 1.325 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 1.985 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445400 ;
    PORT
      LAYER li1 ;
        RECT 1.160 2.030 1.345 2.435 ;
        RECT 1.160 1.855 1.875 2.030 ;
        RECT 1.485 0.825 1.875 1.855 ;
        RECT 1.140 0.655 1.875 0.825 ;
        RECT 1.140 0.255 1.345 0.655 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.085 1.665 0.355 2.435 ;
        RECT 0.525 1.855 0.905 2.635 ;
        RECT 1.515 2.210 1.900 2.635 ;
        RECT 0.085 1.495 1.315 1.665 ;
        RECT 0.085 0.585 0.255 1.495 ;
        RECT 1.015 0.995 1.315 1.495 ;
        RECT 0.085 0.255 0.345 0.585 ;
        RECT 0.605 0.085 0.880 0.565 ;
        RECT 1.515 0.085 1.900 0.485 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkbuf_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__clkbuf_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__clkbuf_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.243000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.755 0.825 1.325 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.995 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.898200 ;
    PORT
      LAYER li1 ;
        RECT 1.145 2.005 1.405 2.465 ;
        RECT 2.105 2.005 2.365 2.465 ;
        RECT 1.145 1.835 2.365 2.005 ;
        RECT 2.105 1.650 2.365 1.835 ;
        RECT 2.105 1.415 2.910 1.650 ;
        RECT 2.410 0.905 2.910 1.415 ;
        RECT 1.050 0.735 2.910 0.905 ;
        RECT 1.050 0.345 1.405 0.735 ;
        RECT 2.105 0.345 2.365 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.085 1.665 0.395 2.465 ;
        RECT 0.615 1.835 0.925 2.635 ;
        RECT 1.625 2.175 1.880 2.635 ;
        RECT 2.545 1.845 2.875 2.635 ;
        RECT 0.085 1.495 1.215 1.665 ;
        RECT 0.085 0.585 0.255 1.495 ;
        RECT 0.995 1.245 1.215 1.495 ;
        RECT 0.995 1.075 2.240 1.245 ;
        RECT 0.085 0.255 0.385 0.585 ;
        RECT 0.605 0.085 0.880 0.565 ;
        RECT 1.625 0.085 1.880 0.565 ;
        RECT 2.585 0.085 2.865 0.565 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkbuf_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__clkbuf_6
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__clkbuf_6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.486000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.715 0.395 1.325 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.275 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.212300 ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.665 1.835 2.460 ;
        RECT 2.445 1.665 2.775 2.460 ;
        RECT 3.385 1.665 3.715 2.460 ;
        RECT 1.505 1.495 4.075 1.665 ;
        RECT 3.745 0.905 4.075 1.495 ;
        RECT 1.505 0.735 4.075 0.905 ;
        RECT 1.505 0.255 1.835 0.735 ;
        RECT 2.445 0.255 2.775 0.735 ;
        RECT 3.385 0.255 3.715 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.095 1.495 0.395 2.635 ;
        RECT 0.565 1.325 0.895 2.465 ;
        RECT 1.065 1.495 1.335 2.635 ;
        RECT 2.005 1.835 2.275 2.635 ;
        RECT 2.945 1.835 3.215 2.635 ;
        RECT 3.885 1.835 4.155 2.635 ;
        RECT 0.565 1.075 3.390 1.325 ;
        RECT 0.145 0.085 0.395 0.545 ;
        RECT 0.565 0.265 0.895 1.075 ;
        RECT 1.065 0.085 1.335 0.610 ;
        RECT 2.005 0.085 2.275 0.565 ;
        RECT 2.945 0.085 3.215 0.565 ;
        RECT 3.885 0.085 4.155 0.565 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkbuf_6

#--------EOF---------

MACRO sky130_fd_sc_hdll__clkbuf_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__clkbuf_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.486000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.715 0.400 1.325 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.320 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.775400 ;
    PORT
      LAYER li1 ;
        RECT 1.570 1.735 1.830 2.460 ;
        RECT 2.530 1.735 2.790 2.460 ;
        RECT 3.490 1.735 3.750 2.460 ;
        RECT 4.450 1.735 4.710 2.460 ;
        RECT 1.570 1.495 5.230 1.735 ;
        RECT 4.160 0.905 5.230 1.495 ;
        RECT 1.570 0.735 5.230 0.905 ;
        RECT 1.570 0.280 1.830 0.735 ;
        RECT 2.530 0.280 2.790 0.735 ;
        RECT 3.490 0.280 3.750 0.735 ;
        RECT 4.450 0.280 4.710 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.095 1.525 0.390 2.635 ;
        RECT 0.620 1.325 0.870 2.460 ;
        RECT 1.090 1.525 1.350 2.635 ;
        RECT 2.050 1.905 2.310 2.635 ;
        RECT 3.010 1.905 3.270 2.635 ;
        RECT 3.970 1.905 4.230 2.635 ;
        RECT 4.930 1.905 5.225 2.635 ;
        RECT 0.620 1.075 3.990 1.325 ;
        RECT 0.145 0.085 0.390 0.545 ;
        RECT 0.620 0.265 0.870 1.075 ;
        RECT 1.090 0.085 1.350 0.610 ;
        RECT 2.050 0.085 2.310 0.565 ;
        RECT 3.010 0.085 3.270 0.565 ;
        RECT 3.970 0.085 4.230 0.565 ;
        RECT 4.930 0.085 5.230 0.565 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkbuf_8

#--------EOF---------

MACRO sky130_fd_sc_hdll__clkbuf_12
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__clkbuf_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.280 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.972000 ;
    PORT
      LAYER li1 ;
        RECT 0.525 1.075 1.320 1.305 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.280 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 8.035 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.470 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.280 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.420400 ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.665 2.745 2.465 ;
        RECT 3.415 1.665 3.685 2.465 ;
        RECT 4.355 1.665 4.625 2.465 ;
        RECT 5.295 1.665 5.565 2.465 ;
        RECT 6.235 1.665 6.505 2.465 ;
        RECT 7.175 1.665 7.445 2.465 ;
        RECT 2.445 1.475 7.445 1.665 ;
        RECT 6.960 0.905 7.445 1.475 ;
        RECT 2.475 0.715 7.445 0.905 ;
        RECT 2.475 0.280 2.745 0.715 ;
        RECT 3.415 0.280 3.685 0.715 ;
        RECT 4.355 0.280 4.625 0.715 ;
        RECT 5.295 0.280 5.565 0.715 ;
        RECT 6.235 0.280 6.505 0.715 ;
        RECT 7.175 0.280 7.445 0.715 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.280 2.805 ;
        RECT 0.095 1.495 0.395 2.635 ;
        RECT 0.565 1.665 0.895 2.465 ;
        RECT 1.065 1.835 1.335 2.635 ;
        RECT 1.535 1.665 1.805 2.465 ;
        RECT 0.565 1.495 1.805 1.665 ;
        RECT 0.570 1.475 1.805 1.495 ;
        RECT 1.975 1.475 2.275 2.635 ;
        RECT 2.915 1.835 3.245 2.635 ;
        RECT 3.855 1.835 4.185 2.635 ;
        RECT 4.795 1.835 5.125 2.635 ;
        RECT 5.735 1.835 6.065 2.635 ;
        RECT 6.675 1.835 7.005 2.635 ;
        RECT 1.535 1.305 1.805 1.475 ;
        RECT 7.615 1.465 7.945 2.635 ;
        RECT 1.535 1.075 6.685 1.305 ;
        RECT 1.535 0.905 1.805 1.075 ;
        RECT 0.595 0.715 1.805 0.905 ;
        RECT 0.095 0.085 0.425 0.610 ;
        RECT 0.595 0.280 0.865 0.715 ;
        RECT 1.035 0.085 1.365 0.545 ;
        RECT 1.535 0.280 1.805 0.715 ;
        RECT 1.975 0.085 2.305 0.545 ;
        RECT 2.915 0.085 3.245 0.545 ;
        RECT 3.855 0.085 4.185 0.545 ;
        RECT 4.795 0.085 5.125 0.545 ;
        RECT 5.735 0.085 6.065 0.545 ;
        RECT 6.675 0.085 7.005 0.545 ;
        RECT 7.615 0.085 7.945 0.610 ;
        RECT 0.000 -0.085 8.280 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkbuf_12

#--------EOF---------

MACRO sky130_fd_sc_hdll__clkbuf_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__clkbuf_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.120 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.972000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.400 1.325 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.120 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 10.110 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.310 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.120 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.529800 ;
    PORT
      LAYER li1 ;
        RECT 2.530 1.735 2.790 2.460 ;
        RECT 3.490 1.735 3.750 2.460 ;
        RECT 4.450 1.735 4.710 2.460 ;
        RECT 5.410 1.735 5.670 2.460 ;
        RECT 6.355 1.735 6.615 2.460 ;
        RECT 7.315 1.735 7.575 2.460 ;
        RECT 8.275 1.735 8.535 2.460 ;
        RECT 2.530 1.720 8.535 1.735 ;
        RECT 9.245 1.720 9.535 2.460 ;
        RECT 2.530 1.495 10.025 1.720 ;
        RECT 8.760 0.905 10.025 1.495 ;
        RECT 2.530 0.735 10.025 0.905 ;
        RECT 2.530 0.280 2.790 0.735 ;
        RECT 3.490 0.280 3.750 0.735 ;
        RECT 4.450 0.280 4.710 0.735 ;
        RECT 5.345 0.280 5.670 0.735 ;
        RECT 6.355 0.280 6.615 0.735 ;
        RECT 7.315 0.280 7.575 0.735 ;
        RECT 8.275 0.280 8.535 0.735 ;
        RECT 9.245 0.280 9.505 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.120 2.805 ;
        RECT 0.095 1.825 0.390 2.635 ;
        RECT 0.620 1.325 0.865 2.465 ;
        RECT 1.090 1.825 1.350 2.635 ;
        RECT 2.050 2.630 9.025 2.635 ;
        RECT 1.580 1.325 1.830 2.460 ;
        RECT 2.050 1.835 2.310 2.630 ;
        RECT 3.010 1.905 3.270 2.630 ;
        RECT 3.970 1.905 4.230 2.630 ;
        RECT 4.930 1.905 5.190 2.630 ;
        RECT 5.890 1.905 6.135 2.630 ;
        RECT 6.850 1.905 7.095 2.630 ;
        RECT 7.810 1.905 8.055 2.630 ;
        RECT 8.770 1.905 9.025 2.630 ;
        RECT 9.755 1.890 10.025 2.635 ;
        RECT 0.620 1.075 8.540 1.325 ;
        RECT 0.085 0.085 0.390 0.595 ;
        RECT 0.620 0.265 0.870 1.075 ;
        RECT 1.090 0.085 1.350 0.610 ;
        RECT 1.580 0.265 1.830 1.075 ;
        RECT 2.050 0.085 2.310 0.645 ;
        RECT 3.010 0.085 3.270 0.565 ;
        RECT 3.970 0.085 4.230 0.565 ;
        RECT 4.930 0.085 5.175 0.565 ;
        RECT 5.890 0.085 6.135 0.565 ;
        RECT 6.845 0.085 7.095 0.565 ;
        RECT 7.805 0.085 8.055 0.565 ;
        RECT 8.765 0.085 9.025 0.565 ;
        RECT 9.725 0.085 10.025 0.565 ;
        RECT 0.000 -0.085 10.120 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkbuf_16

#--------EOF---------

MACRO sky130_fd_sc_hdll__clkinv_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__clkinv_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.375 0.325 1.325 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.375900 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.290 0.895 2.465 ;
        RECT 0.515 0.760 1.395 1.290 ;
        RECT 0.515 0.255 0.890 0.760 ;
    END
  END Y
  OBS
      LAYER pwell ;
        RECT 0.470 0.105 1.480 0.785 ;
      LAYER li1 ;
        RECT 0.000 2.635 1.840 2.805 ;
        RECT 0.085 1.665 0.345 2.635 ;
        RECT 1.115 1.665 1.395 2.635 ;
        RECT 1.115 0.085 1.395 0.590 ;
        RECT 0.000 -0.085 1.840 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkinv_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__clkinv_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__clkinv_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.065 1.335 1.290 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.728600 ;
    PORT
      LAYER li1 ;
        RECT 0.155 1.630 0.410 2.435 ;
        RECT 1.110 1.630 1.370 2.435 ;
        RECT 0.155 1.460 2.155 1.630 ;
        RECT 1.520 0.895 2.155 1.460 ;
        RECT 1.125 0.725 2.155 0.895 ;
        RECT 1.125 0.280 1.350 0.725 ;
    END
  END Y
  OBS
      LAYER pwell ;
        RECT 0.520 0.105 1.985 0.785 ;
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.630 1.800 0.890 2.635 ;
        RECT 1.605 1.800 1.860 2.635 ;
        RECT 0.560 0.085 0.905 0.610 ;
        RECT 1.520 0.085 1.900 0.555 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkinv_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__clkinv_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__clkinv_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332000 ;
    PORT
      LAYER li1 ;
        RECT 0.445 1.065 2.910 1.290 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.177200 ;
    PORT
      LAYER li1 ;
        RECT 0.655 1.630 0.910 2.435 ;
        RECT 1.615 1.630 1.870 2.435 ;
        RECT 2.570 1.630 2.830 2.435 ;
        RECT 0.105 1.460 3.570 1.630 ;
        RECT 0.105 0.895 0.275 1.460 ;
        RECT 3.270 0.895 3.570 1.460 ;
        RECT 0.105 0.725 3.570 0.895 ;
        RECT 1.130 0.280 1.390 0.725 ;
        RECT 2.090 0.280 2.345 0.725 ;
    END
  END Y
  OBS
      LAYER pwell ;
        RECT 0.410 0.105 3.085 0.785 ;
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.085 1.800 0.430 2.635 ;
        RECT 1.130 1.800 1.390 2.635 ;
        RECT 2.090 1.800 2.350 2.635 ;
        RECT 3.050 1.800 3.435 2.635 ;
        RECT 0.565 0.085 0.910 0.555 ;
        RECT 1.610 0.085 1.870 0.555 ;
        RECT 2.565 0.085 2.865 0.555 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkinv_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__clkinv_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__clkinv_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.664000 ;
    PORT
      LAYER li1 ;
        RECT 0.455 1.035 5.565 1.290 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150 -0.085 0.320 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.386400 ;
    PORT
      LAYER li1 ;
        RECT 0.615 1.630 0.855 2.435 ;
        RECT 1.555 1.630 1.795 2.435 ;
        RECT 2.495 1.630 2.745 2.435 ;
        RECT 3.430 1.630 3.675 2.435 ;
        RECT 4.420 1.630 4.725 2.435 ;
        RECT 5.465 1.630 5.705 2.435 ;
        RECT 0.115 1.460 6.330 1.630 ;
        RECT 0.115 0.865 0.285 1.460 ;
        RECT 6.060 0.865 6.330 1.460 ;
        RECT 0.115 0.695 6.330 0.865 ;
        RECT 1.685 0.280 1.875 0.695 ;
        RECT 2.645 0.280 2.835 0.695 ;
        RECT 3.605 0.280 3.795 0.695 ;
        RECT 4.665 0.280 4.855 0.695 ;
    END
  END Y
  OBS
      LAYER pwell ;
        RECT 1.045 0.105 5.595 0.785 ;
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.135 1.800 0.395 2.635 ;
        RECT 1.075 1.800 1.335 2.635 ;
        RECT 2.015 1.800 2.275 2.635 ;
        RECT 2.965 1.800 3.210 2.635 ;
        RECT 3.895 1.800 4.200 2.635 ;
        RECT 4.945 1.800 5.245 2.635 ;
        RECT 5.925 1.800 6.180 2.635 ;
        RECT 1.135 0.085 1.465 0.525 ;
        RECT 2.095 0.085 2.425 0.525 ;
        RECT 3.055 0.085 3.435 0.525 ;
        RECT 4.015 0.085 4.445 0.525 ;
        RECT 5.075 0.085 5.505 0.525 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkinv_8

#--------EOF---------

MACRO sky130_fd_sc_hdll__clkinv_12
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__clkinv_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.200 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.996000 ;
    PORT
      LAYER li1 ;
        RECT 0.455 1.035 7.925 1.290 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.200 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150 -0.085 0.320 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.390 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.200 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.290400 ;
    PORT
      LAYER li1 ;
        RECT 0.595 1.630 0.865 2.465 ;
        RECT 1.535 1.630 1.805 2.465 ;
        RECT 2.475 1.630 2.745 2.465 ;
        RECT 3.415 1.630 3.685 2.465 ;
        RECT 4.355 1.630 4.625 2.465 ;
        RECT 5.295 1.630 5.565 2.465 ;
        RECT 6.235 1.630 6.505 2.465 ;
        RECT 7.175 1.630 7.445 2.465 ;
        RECT 8.115 1.630 8.385 2.465 ;
        RECT 0.115 1.460 8.655 1.630 ;
        RECT 0.115 0.865 0.285 1.460 ;
        RECT 8.100 0.865 8.655 1.460 ;
        RECT 0.115 0.695 8.655 0.865 ;
        RECT 2.005 0.255 2.275 0.695 ;
        RECT 2.945 0.255 3.215 0.695 ;
        RECT 3.885 0.255 4.155 0.695 ;
        RECT 4.825 0.255 5.095 0.695 ;
        RECT 5.765 0.255 6.035 0.695 ;
        RECT 6.705 0.255 6.975 0.695 ;
    END
  END Y
  OBS
      LAYER pwell ;
        RECT 1.075 0.105 7.905 0.785 ;
      LAYER li1 ;
        RECT 0.000 2.635 9.200 2.805 ;
        RECT 0.095 1.800 0.425 2.635 ;
        RECT 1.035 1.800 1.365 2.635 ;
        RECT 1.975 1.800 2.305 2.635 ;
        RECT 2.915 1.800 3.245 2.635 ;
        RECT 3.855 1.800 4.185 2.635 ;
        RECT 4.795 1.800 5.125 2.635 ;
        RECT 5.735 1.800 6.065 2.635 ;
        RECT 6.675 1.800 7.005 2.635 ;
        RECT 7.615 1.800 7.945 2.635 ;
        RECT 8.555 1.800 8.885 2.635 ;
        RECT 1.165 0.085 1.835 0.525 ;
        RECT 2.445 0.085 2.775 0.525 ;
        RECT 3.385 0.085 3.715 0.525 ;
        RECT 4.325 0.085 4.655 0.525 ;
        RECT 5.265 0.085 5.595 0.525 ;
        RECT 6.205 0.085 6.535 0.525 ;
        RECT 7.145 0.085 7.815 0.525 ;
        RECT 0.000 -0.085 9.200 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkinv_12

#--------EOF---------

MACRO sky130_fd_sc_hdll__clkinv_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__clkinv_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.420 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.328000 ;
    PORT
      LAYER met1 ;
        RECT 1.615 1.260 2.415 1.305 ;
        RECT 10.285 1.260 11.135 1.305 ;
        RECT 1.615 1.120 11.135 1.260 ;
        RECT 1.615 1.075 2.415 1.120 ;
        RECT 10.285 1.075 11.135 1.120 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 12.420 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 12.610 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 12.420 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.928900 ;
    PORT
      LAYER li1 ;
        RECT 0.625 1.665 0.880 2.465 ;
        RECT 1.585 1.665 1.840 2.450 ;
        RECT 2.575 1.665 2.800 2.465 ;
        RECT 3.505 1.665 3.760 2.450 ;
        RECT 4.465 1.665 4.705 2.450 ;
        RECT 5.455 1.665 5.830 2.450 ;
        RECT 6.575 1.665 6.825 2.450 ;
        RECT 7.535 1.665 7.785 2.450 ;
        RECT 8.495 1.665 8.745 2.450 ;
        RECT 9.455 1.665 9.705 2.450 ;
        RECT 10.415 1.665 10.655 2.450 ;
        RECT 11.375 1.665 11.630 2.450 ;
        RECT 0.625 1.455 11.630 1.665 ;
        RECT 2.575 1.415 9.705 1.455 ;
        RECT 2.575 0.280 2.800 1.415 ;
        RECT 3.505 0.280 3.760 1.415 ;
        RECT 4.465 0.280 4.705 1.415 ;
        RECT 5.455 0.280 5.805 1.415 ;
        RECT 6.575 0.280 6.825 1.415 ;
        RECT 7.535 0.280 7.785 1.415 ;
        RECT 8.495 0.280 8.745 1.415 ;
        RECT 9.455 0.280 9.705 1.415 ;
    END
  END Y
  OBS
      LAYER pwell ;
        RECT 1.935 0.105 10.315 0.785 ;
      LAYER li1 ;
        RECT 0.000 2.635 12.420 2.805 ;
        RECT 0.140 1.495 0.405 2.635 ;
        RECT 1.100 1.835 1.360 2.635 ;
        RECT 2.065 1.835 2.320 2.635 ;
        RECT 3.020 1.835 3.280 2.635 ;
        RECT 3.985 1.835 4.240 2.635 ;
        RECT 4.965 1.835 5.220 2.635 ;
        RECT 6.090 2.120 6.350 2.635 ;
        RECT 6.090 1.835 6.345 2.120 ;
        RECT 7.055 1.835 7.310 2.635 ;
        RECT 8.015 1.835 8.270 2.635 ;
        RECT 8.975 1.835 9.230 2.635 ;
        RECT 9.935 1.835 10.190 2.635 ;
        RECT 10.895 1.835 11.150 2.635 ;
        RECT 11.850 1.835 12.110 2.635 ;
        RECT 0.345 0.895 2.355 1.275 ;
        RECT 9.930 0.895 11.910 1.275 ;
        RECT 2.055 0.085 2.325 0.610 ;
        RECT 3.020 0.085 3.285 0.610 ;
        RECT 3.980 0.085 4.245 0.610 ;
        RECT 4.965 0.085 5.230 0.610 ;
        RECT 6.090 0.085 6.355 0.610 ;
        RECT 7.050 0.085 7.275 0.610 ;
        RECT 8.010 0.085 8.275 0.610 ;
        RECT 8.970 0.085 9.235 0.610 ;
        RECT 9.930 0.085 10.195 0.610 ;
        RECT 0.000 -0.085 12.420 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 1.675 1.105 1.845 1.275 ;
        RECT 2.185 1.105 2.355 1.275 ;
        RECT 10.395 1.105 10.565 1.275 ;
        RECT 10.905 1.105 11.075 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkinv_16

#--------EOF---------

MACRO sky130_fd_sc_hdll__clkinvlp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__clkinvlp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.665000 ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.995 0.600 1.665 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.185 0.205 1.675 1.015 ;
        RECT 0.185 0.085 0.315 0.205 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.436750 ;
    PORT
      LAYER li1 ;
        RECT 0.785 0.750 1.235 2.455 ;
        RECT 0.785 0.315 1.545 0.750 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.840 2.805 ;
        RECT 0.225 2.625 1.665 2.635 ;
        RECT 0.225 1.835 0.555 2.625 ;
        RECT 1.405 1.455 1.665 2.625 ;
        RECT 0.295 0.085 0.615 0.745 ;
        RECT 0.000 -0.085 1.840 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkinvlp_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__clkinvlp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__clkinvlp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.330000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.745 0.425 1.325 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.090 0.915 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.694000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.295 0.945 2.465 ;
        RECT 1.655 1.295 1.985 2.465 ;
        RECT 0.605 1.015 1.985 1.295 ;
        RECT 0.605 0.680 0.955 1.015 ;
        RECT 0.605 0.255 1.165 0.680 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.095 1.495 0.420 2.635 ;
        RECT 1.185 1.465 1.460 2.635 ;
        RECT 2.225 1.465 2.505 2.635 ;
        RECT 0.095 0.085 0.425 0.575 ;
        RECT 1.675 0.085 2.000 0.775 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkinvlp_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__clkmux2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__clkmux2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.232200 ;
    PORT
      LAYER li1 ;
        RECT 2.290 0.255 2.615 1.415 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.232200 ;
    PORT
      LAYER li1 ;
        RECT 1.780 1.615 3.075 1.785 ;
        RECT 1.780 0.810 1.950 1.615 ;
        RECT 2.785 0.255 3.075 1.615 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.479400 ;
    PORT
      LAYER li1 ;
        RECT 1.070 2.295 3.415 2.465 ;
        RECT 1.070 1.325 1.270 2.295 ;
        RECT 3.245 1.630 3.415 2.295 ;
        RECT 3.245 1.440 3.995 1.630 ;
        RECT 0.995 0.995 1.270 1.325 ;
        RECT 3.805 1.055 3.995 1.440 ;
    END
  END S
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.785 0.985 0.885 ;
        RECT 3.485 0.785 4.405 0.885 ;
        RECT 0.005 0.105 4.405 0.785 ;
        RECT 0.420 -0.085 0.640 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.405200 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.495 0.425 2.465 ;
        RECT 0.090 0.255 0.345 1.495 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.645 1.495 0.815 2.635 ;
        RECT 1.440 1.955 2.885 2.125 ;
        RECT 0.515 0.825 0.685 1.325 ;
        RECT 1.440 0.825 1.610 1.955 ;
        RECT 3.585 1.835 3.815 2.635 ;
        RECT 3.985 1.835 4.385 2.465 ;
        RECT 0.515 0.655 1.610 0.825 ;
        RECT 3.325 0.865 3.495 1.185 ;
        RECT 4.215 0.865 4.385 1.835 ;
        RECT 3.325 0.695 4.385 0.865 ;
        RECT 1.435 0.620 1.610 0.655 ;
        RECT 0.515 0.085 0.895 0.485 ;
        RECT 1.435 0.255 1.955 0.620 ;
        RECT 3.250 0.085 3.765 0.525 ;
        RECT 4.035 0.255 4.280 0.695 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkmux2_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__clkmux2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__clkmux2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.232200 ;
    PORT
      LAYER li1 ;
        RECT 2.750 0.255 3.075 1.415 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.232200 ;
    PORT
      LAYER li1 ;
        RECT 2.240 1.615 3.535 1.785 ;
        RECT 2.240 0.810 2.410 1.615 ;
        RECT 3.245 0.255 3.535 1.615 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.479400 ;
    PORT
      LAYER li1 ;
        RECT 1.530 2.295 3.875 2.465 ;
        RECT 1.530 1.325 1.730 2.295 ;
        RECT 3.705 1.630 3.875 2.295 ;
        RECT 3.705 1.440 4.455 1.630 ;
        RECT 1.455 0.995 1.730 1.325 ;
        RECT 4.265 1.055 4.455 1.440 ;
    END
  END S
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.785 1.445 0.885 ;
        RECT 3.945 0.785 4.865 0.885 ;
        RECT 0.005 0.105 4.865 0.785 ;
        RECT 0.880 -0.085 1.100 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.430400 ;
    PORT
      LAYER li1 ;
        RECT 0.555 1.495 0.895 2.465 ;
        RECT 0.555 0.255 0.805 1.495 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.060 2.805 ;
        RECT 0.135 1.495 0.380 2.635 ;
        RECT 1.075 1.495 1.325 2.635 ;
        RECT 1.900 1.955 3.345 2.125 ;
        RECT 0.975 0.825 1.145 1.325 ;
        RECT 1.900 0.825 2.070 1.955 ;
        RECT 4.045 1.835 4.275 2.635 ;
        RECT 4.445 1.835 4.845 2.465 ;
        RECT 0.975 0.655 2.070 0.825 ;
        RECT 3.785 0.865 3.955 1.185 ;
        RECT 4.675 0.865 4.845 1.835 ;
        RECT 3.785 0.695 4.845 0.865 ;
        RECT 0.135 0.085 0.385 0.655 ;
        RECT 1.895 0.620 2.070 0.655 ;
        RECT 0.975 0.085 1.355 0.485 ;
        RECT 1.895 0.255 2.580 0.620 ;
        RECT 3.710 0.085 4.225 0.525 ;
        RECT 4.495 0.255 4.740 0.695 ;
        RECT 0.000 -0.085 5.060 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkmux2_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__clkmux2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__clkmux2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.232200 ;
    PORT
      LAYER li1 ;
        RECT 3.670 0.255 3.995 1.415 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.232200 ;
    PORT
      LAYER li1 ;
        RECT 3.160 1.615 4.455 1.785 ;
        RECT 3.160 0.810 3.330 1.615 ;
        RECT 4.165 0.255 4.455 1.615 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.479400 ;
    PORT
      LAYER li1 ;
        RECT 2.450 2.295 4.795 2.465 ;
        RECT 2.450 1.325 2.650 2.295 ;
        RECT 4.625 1.630 4.795 2.295 ;
        RECT 4.625 1.440 5.375 1.630 ;
        RECT 2.375 0.995 2.650 1.325 ;
        RECT 5.185 1.055 5.375 1.440 ;
    END
  END S
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.045 0.785 2.365 0.885 ;
        RECT 4.865 0.785 5.785 0.885 ;
        RECT 0.045 0.105 5.785 0.785 ;
        RECT 1.800 -0.085 2.020 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.860800 ;
    PORT
      LAYER li1 ;
        RECT 0.565 1.495 0.895 2.465 ;
        RECT 1.475 1.495 1.835 2.465 ;
        RECT 0.590 1.325 0.850 1.495 ;
        RECT 1.475 1.325 1.745 1.495 ;
        RECT 0.590 1.065 1.745 1.325 ;
        RECT 0.590 0.255 0.850 1.065 ;
        RECT 1.475 0.255 1.745 1.065 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.135 1.495 0.395 2.635 ;
        RECT 1.065 1.495 1.305 2.635 ;
        RECT 2.005 1.495 2.280 2.635 ;
        RECT 2.820 1.955 4.265 2.125 ;
        RECT 1.915 0.825 2.085 1.325 ;
        RECT 2.820 0.825 2.990 1.955 ;
        RECT 4.965 1.835 5.195 2.635 ;
        RECT 5.365 1.835 5.765 2.465 ;
        RECT 1.915 0.655 2.990 0.825 ;
        RECT 4.705 0.865 4.875 1.185 ;
        RECT 5.595 0.865 5.765 1.835 ;
        RECT 4.705 0.695 5.765 0.865 ;
        RECT 0.175 0.085 0.420 0.655 ;
        RECT 1.055 0.085 1.305 0.655 ;
        RECT 2.815 0.620 2.990 0.655 ;
        RECT 1.915 0.085 2.275 0.485 ;
        RECT 2.815 0.255 3.500 0.620 ;
        RECT 4.630 0.085 5.145 0.525 ;
        RECT 5.415 0.255 5.660 0.695 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkmux2_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__conb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__conb_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 1.570 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  PIN HI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.605 1.740 ;
    END
  END HI
  PIN LO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.775 0.915 1.295 2.465 ;
    END
  END LO
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.380 2.805 ;
        RECT 0.275 1.910 0.605 2.635 ;
        RECT 0.775 0.085 1.115 0.745 ;
        RECT 0.000 -0.085 1.380 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__conb_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__decap_3
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hdll__decap_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 1.375 0.915 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 1.570 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.380 2.805 ;
        RECT 0.085 1.545 1.295 2.635 ;
        RECT 0.085 0.835 0.605 1.375 ;
        RECT 0.775 1.005 1.295 1.545 ;
        RECT 0.085 0.085 1.295 0.835 ;
        RECT 0.000 -0.085 1.380 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__decap_3

#--------EOF---------

MACRO sky130_fd_sc_hdll__decap_4
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hdll__decap_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 1.835 0.915 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.840 2.805 ;
        RECT 0.085 1.545 1.755 2.635 ;
        RECT 0.085 0.855 0.835 1.375 ;
        RECT 1.005 1.025 1.755 1.545 ;
        RECT 0.085 0.085 1.755 0.855 ;
        RECT 0.000 -0.085 1.840 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__decap_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__decap_6
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hdll__decap_6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.755 0.915 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.085 1.545 2.675 2.635 ;
        RECT 0.085 0.855 1.295 1.375 ;
        RECT 1.465 1.025 2.675 1.545 ;
        RECT 0.085 0.085 2.675 0.855 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__decap_6

#--------EOF---------

MACRO sky130_fd_sc_hdll__decap_8
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hdll__decap_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.675 0.915 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.085 1.545 3.595 2.635 ;
        RECT 0.085 0.855 1.735 1.375 ;
        RECT 1.905 1.025 3.595 1.545 ;
        RECT 0.085 0.085 3.595 0.855 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__decap_8

#--------EOF---------

MACRO sky130_fd_sc_hdll__decap_12
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hdll__decap_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.515 0.915 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.085 1.545 5.430 2.635 ;
        RECT 0.085 0.855 2.665 1.375 ;
        RECT 2.835 1.025 5.430 1.545 ;
        RECT 0.085 0.085 5.430 0.855 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__decap_12

#--------EOF---------

MACRO sky130_fd_sc_hdll__dfrtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__dfrtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.660 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.975 0.440 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.455 1.665 1.770 2.005 ;
        RECT 1.455 0.615 1.905 1.665 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277200 ;
    PORT
      LAYER met1 ;
        RECT 3.995 0.920 4.745 0.965 ;
        RECT 7.575 0.920 7.865 0.965 ;
        RECT 3.995 0.780 7.865 0.920 ;
        RECT 3.995 0.735 4.745 0.780 ;
        RECT 7.575 0.735 7.865 0.780 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.660 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.565 0.785 5.545 1.005 ;
        RECT 8.640 0.785 9.640 1.015 ;
        RECT 0.005 0.105 9.640 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.850 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.660 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.472000 ;
    PORT
      LAYER li1 ;
        RECT 9.240 0.255 9.575 2.465 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.660 2.805 ;
        RECT 0.090 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.895 2.635 ;
        RECT 0.090 1.795 0.890 1.965 ;
        RECT 0.660 0.805 0.890 1.795 ;
        RECT 0.090 0.635 0.890 0.805 ;
        RECT 0.090 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.115 0.345 1.285 2.465 ;
        RECT 1.770 2.175 1.940 2.635 ;
        RECT 2.170 2.135 2.420 2.465 ;
        RECT 2.685 2.135 3.365 2.465 ;
        RECT 2.170 2.005 2.340 2.135 ;
        RECT 2.075 1.835 2.340 2.005 ;
        RECT 2.075 0.475 2.245 1.835 ;
        RECT 2.510 1.575 3.025 1.965 ;
        RECT 2.425 0.765 2.685 1.385 ;
        RECT 2.855 0.985 3.025 1.575 ;
        RECT 3.195 1.355 3.365 2.135 ;
        RECT 3.535 2.035 3.705 2.375 ;
        RECT 3.990 2.205 4.320 2.635 ;
        RECT 4.540 2.035 4.710 2.375 ;
        RECT 5.005 2.175 5.425 2.635 ;
        RECT 3.535 1.865 4.710 2.035 ;
        RECT 5.645 2.005 5.815 2.465 ;
        RECT 6.050 2.125 7.005 2.465 ;
        RECT 7.340 2.175 7.590 2.635 ;
        RECT 5.155 1.835 5.815 2.005 ;
        RECT 5.155 1.695 5.325 1.835 ;
        RECT 3.725 1.525 5.325 1.695 ;
        RECT 6.145 1.665 6.660 1.955 ;
        RECT 3.195 1.185 4.985 1.355 ;
        RECT 2.855 0.765 3.210 0.985 ;
        RECT 3.430 0.475 3.600 1.185 ;
        RECT 3.805 0.765 4.645 1.015 ;
        RECT 4.815 1.005 4.985 1.185 ;
        RECT 5.155 0.835 5.325 1.525 ;
        RECT 1.575 0.085 1.905 0.445 ;
        RECT 2.075 0.305 2.495 0.475 ;
        RECT 2.695 0.305 3.600 0.475 ;
        RECT 4.525 0.085 4.855 0.545 ;
        RECT 5.065 0.445 5.325 0.835 ;
        RECT 5.605 1.655 6.660 1.665 ;
        RECT 6.835 1.745 7.005 2.125 ;
        RECT 7.810 2.085 7.980 2.375 ;
        RECT 8.160 2.255 8.540 2.635 ;
        RECT 7.810 1.915 8.610 2.085 ;
        RECT 5.605 1.495 6.315 1.655 ;
        RECT 6.835 1.575 8.270 1.745 ;
        RECT 5.605 0.705 5.775 1.495 ;
        RECT 6.835 1.485 7.055 1.575 ;
        RECT 5.945 0.705 6.315 1.325 ;
        RECT 6.485 1.315 7.055 1.485 ;
        RECT 6.485 0.535 6.655 1.315 ;
        RECT 6.955 0.865 7.225 1.145 ;
        RECT 6.955 0.695 7.335 0.865 ;
        RECT 5.065 0.275 5.465 0.445 ;
        RECT 5.735 0.255 6.655 0.535 ;
        RECT 6.825 0.085 6.995 0.525 ;
        RECT 7.165 0.465 7.335 0.695 ;
        RECT 7.505 0.635 7.905 1.405 ;
        RECT 8.440 1.295 8.610 1.915 ;
        RECT 8.810 1.575 8.980 2.635 ;
        RECT 8.290 1.285 8.610 1.295 ;
        RECT 8.290 1.075 9.070 1.285 ;
        RECT 8.290 0.465 8.635 1.075 ;
        RECT 7.165 0.295 8.635 0.465 ;
        RECT 8.810 0.085 8.980 0.895 ;
        RECT 0.000 -0.085 9.660 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 0.660 1.105 0.830 1.275 ;
        RECT 1.115 1.785 1.285 1.955 ;
        RECT 2.725 1.785 2.895 1.955 ;
        RECT 2.480 1.105 2.650 1.275 ;
        RECT 6.470 1.785 6.640 1.955 ;
        RECT 4.105 0.765 4.275 0.935 ;
        RECT 4.465 0.765 4.635 0.935 ;
        RECT 6.020 1.105 6.190 1.275 ;
        RECT 7.635 0.765 7.805 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
      LAYER met1 ;
        RECT 1.005 1.940 1.345 1.985 ;
        RECT 2.665 1.940 2.955 1.985 ;
        RECT 6.410 1.940 6.700 1.985 ;
        RECT 1.005 1.800 6.700 1.940 ;
        RECT 1.005 1.755 1.345 1.800 ;
        RECT 2.665 1.755 2.955 1.800 ;
        RECT 6.410 1.755 6.700 1.800 ;
        RECT 0.600 1.260 0.890 1.305 ;
        RECT 2.420 1.260 2.710 1.305 ;
        RECT 5.960 1.260 6.250 1.305 ;
        RECT 0.600 1.120 6.250 1.260 ;
        RECT 0.600 1.075 0.890 1.120 ;
        RECT 2.420 1.075 2.710 1.120 ;
        RECT 5.960 1.075 6.250 1.120 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dfrtp_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__dfrtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__dfrtp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.120 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.975 0.440 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.455 1.665 1.770 2.005 ;
        RECT 1.455 0.615 1.905 1.665 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277200 ;
    PORT
      LAYER met1 ;
        RECT 3.995 0.920 4.745 0.965 ;
        RECT 7.575 0.920 7.865 0.965 ;
        RECT 3.995 0.780 7.865 0.920 ;
        RECT 3.995 0.735 4.745 0.780 ;
        RECT 7.575 0.735 7.865 0.780 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.120 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.565 0.785 5.545 1.005 ;
        RECT 8.640 0.785 10.090 1.015 ;
        RECT 0.005 0.105 10.090 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.310 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.120 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.530500 ;
    PORT
      LAYER li1 ;
        RECT 9.240 1.625 9.530 2.465 ;
        RECT 9.240 1.455 10.010 1.625 ;
        RECT 9.625 0.905 10.010 1.455 ;
        RECT 9.150 0.735 10.010 0.905 ;
        RECT 9.150 0.255 9.530 0.735 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.120 2.805 ;
        RECT 0.090 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.895 2.635 ;
        RECT 0.090 1.795 0.890 1.965 ;
        RECT 0.660 0.805 0.890 1.795 ;
        RECT 0.090 0.635 0.890 0.805 ;
        RECT 0.090 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.115 0.345 1.285 2.465 ;
        RECT 1.770 2.175 1.940 2.635 ;
        RECT 2.170 2.135 2.420 2.465 ;
        RECT 2.685 2.135 3.365 2.465 ;
        RECT 2.170 2.005 2.340 2.135 ;
        RECT 2.075 1.835 2.340 2.005 ;
        RECT 2.075 0.475 2.245 1.835 ;
        RECT 2.510 1.575 3.025 1.965 ;
        RECT 2.425 0.765 2.685 1.385 ;
        RECT 2.855 0.985 3.025 1.575 ;
        RECT 3.195 1.355 3.365 2.135 ;
        RECT 3.535 2.035 3.705 2.375 ;
        RECT 3.990 2.205 4.320 2.635 ;
        RECT 4.540 2.035 4.710 2.375 ;
        RECT 5.005 2.175 5.425 2.635 ;
        RECT 3.535 1.865 4.710 2.035 ;
        RECT 5.645 2.005 5.815 2.465 ;
        RECT 6.050 2.125 7.005 2.465 ;
        RECT 7.340 2.175 7.590 2.635 ;
        RECT 5.155 1.835 5.815 2.005 ;
        RECT 5.155 1.695 5.325 1.835 ;
        RECT 3.725 1.525 5.325 1.695 ;
        RECT 6.145 1.665 6.660 1.955 ;
        RECT 3.195 1.185 4.985 1.355 ;
        RECT 2.855 0.765 3.210 0.985 ;
        RECT 3.430 0.475 3.600 1.185 ;
        RECT 3.805 0.765 4.645 1.015 ;
        RECT 4.815 1.005 4.985 1.185 ;
        RECT 5.155 0.835 5.325 1.525 ;
        RECT 1.575 0.085 1.905 0.445 ;
        RECT 2.075 0.305 2.495 0.475 ;
        RECT 2.695 0.305 3.600 0.475 ;
        RECT 4.525 0.085 4.855 0.545 ;
        RECT 5.065 0.445 5.325 0.835 ;
        RECT 5.605 1.655 6.660 1.665 ;
        RECT 6.835 1.745 7.005 2.125 ;
        RECT 7.810 2.085 7.980 2.375 ;
        RECT 8.160 2.255 8.540 2.635 ;
        RECT 7.810 1.915 8.610 2.085 ;
        RECT 5.605 1.495 6.315 1.655 ;
        RECT 6.835 1.575 8.270 1.745 ;
        RECT 5.605 0.705 5.775 1.495 ;
        RECT 6.835 1.485 7.055 1.575 ;
        RECT 5.945 0.705 6.315 1.325 ;
        RECT 6.485 1.315 7.055 1.485 ;
        RECT 6.485 0.535 6.655 1.315 ;
        RECT 6.955 0.865 7.225 1.145 ;
        RECT 6.955 0.695 7.335 0.865 ;
        RECT 5.065 0.275 5.465 0.445 ;
        RECT 5.735 0.255 6.655 0.535 ;
        RECT 6.825 0.085 6.995 0.525 ;
        RECT 7.165 0.465 7.335 0.695 ;
        RECT 7.505 0.635 7.905 1.405 ;
        RECT 8.440 1.295 8.610 1.915 ;
        RECT 8.810 1.575 8.980 2.635 ;
        RECT 9.750 1.795 9.920 2.635 ;
        RECT 8.290 1.285 8.610 1.295 ;
        RECT 8.290 1.075 9.335 1.285 ;
        RECT 8.290 0.465 8.635 1.075 ;
        RECT 7.165 0.295 8.635 0.465 ;
        RECT 8.810 0.085 8.980 0.895 ;
        RECT 9.750 0.085 9.920 0.555 ;
        RECT 0.000 -0.085 10.120 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 0.660 1.105 0.830 1.275 ;
        RECT 1.115 1.785 1.285 1.955 ;
        RECT 2.725 1.785 2.895 1.955 ;
        RECT 2.480 1.105 2.650 1.275 ;
        RECT 6.470 1.785 6.640 1.955 ;
        RECT 4.105 0.765 4.275 0.935 ;
        RECT 4.465 0.765 4.635 0.935 ;
        RECT 6.020 1.105 6.190 1.275 ;
        RECT 7.635 0.765 7.805 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
      LAYER met1 ;
        RECT 1.005 1.940 1.345 1.985 ;
        RECT 2.665 1.940 2.955 1.985 ;
        RECT 6.410 1.940 6.700 1.985 ;
        RECT 1.005 1.800 6.700 1.940 ;
        RECT 1.005 1.755 1.345 1.800 ;
        RECT 2.665 1.755 2.955 1.800 ;
        RECT 6.410 1.755 6.700 1.800 ;
        RECT 0.600 1.260 0.890 1.305 ;
        RECT 2.420 1.260 2.710 1.305 ;
        RECT 5.960 1.260 6.250 1.305 ;
        RECT 0.600 1.120 6.250 1.260 ;
        RECT 0.600 1.075 0.890 1.120 ;
        RECT 2.420 1.075 2.710 1.120 ;
        RECT 5.960 1.075 6.250 1.120 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dfrtp_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__dfrtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__dfrtp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.500 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.975 0.440 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.455 1.665 1.780 2.450 ;
        RECT 1.455 0.615 1.975 1.665 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277200 ;
    PORT
      LAYER met1 ;
        RECT 4.175 0.920 4.925 0.965 ;
        RECT 7.810 0.920 8.395 1.280 ;
        RECT 4.175 0.780 8.395 0.920 ;
        RECT 4.175 0.735 4.925 0.780 ;
        RECT 8.105 0.735 8.395 0.780 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.500 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.865 0.785 5.845 1.005 ;
        RECT 8.965 0.785 11.375 1.015 ;
        RECT 0.005 0.105 11.375 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 11.690 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.500 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.996000 ;
    PORT
      LAYER li1 ;
        RECT 9.565 1.625 9.855 2.465 ;
        RECT 10.505 1.625 10.755 2.465 ;
        RECT 9.565 1.455 11.405 1.625 ;
        RECT 10.995 0.905 11.405 1.455 ;
        RECT 9.475 0.735 11.405 0.905 ;
        RECT 9.475 0.255 9.855 0.735 ;
        RECT 10.415 0.255 10.795 0.735 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 11.500 2.805 ;
        RECT 0.090 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.895 2.635 ;
        RECT 0.090 1.795 0.890 1.965 ;
        RECT 0.660 0.805 0.890 1.795 ;
        RECT 0.090 0.635 0.890 0.805 ;
        RECT 0.090 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.115 0.345 1.285 2.465 ;
        RECT 1.950 2.175 2.200 2.635 ;
        RECT 2.420 2.135 2.670 2.465 ;
        RECT 2.935 2.135 3.665 2.465 ;
        RECT 2.420 2.005 2.590 2.135 ;
        RECT 2.145 1.835 2.590 2.005 ;
        RECT 2.145 0.475 2.315 1.835 ;
        RECT 2.760 1.575 3.275 1.965 ;
        RECT 2.535 0.765 2.935 1.385 ;
        RECT 3.105 0.985 3.275 1.575 ;
        RECT 3.495 1.355 3.665 2.135 ;
        RECT 3.835 2.035 4.005 2.375 ;
        RECT 4.290 2.205 4.620 2.635 ;
        RECT 4.840 2.035 5.010 2.375 ;
        RECT 5.305 2.175 5.725 2.635 ;
        RECT 3.835 1.865 5.010 2.035 ;
        RECT 5.945 2.005 6.115 2.465 ;
        RECT 6.350 2.125 7.470 2.465 ;
        RECT 7.640 2.175 7.890 2.635 ;
        RECT 5.505 1.835 6.115 2.005 ;
        RECT 5.505 1.695 5.675 1.835 ;
        RECT 4.025 1.525 5.675 1.695 ;
        RECT 6.470 1.665 7.030 1.955 ;
        RECT 3.495 1.185 5.285 1.355 ;
        RECT 3.105 0.765 3.510 0.985 ;
        RECT 3.680 0.475 3.850 1.185 ;
        RECT 4.175 0.765 4.945 1.015 ;
        RECT 5.115 1.005 5.285 1.185 ;
        RECT 5.505 0.835 5.675 1.525 ;
        RECT 1.645 0.085 1.975 0.445 ;
        RECT 2.145 0.305 2.690 0.475 ;
        RECT 2.945 0.305 3.850 0.475 ;
        RECT 4.825 0.085 5.155 0.545 ;
        RECT 5.365 0.445 5.675 0.835 ;
        RECT 5.915 1.655 7.030 1.665 ;
        RECT 7.250 1.745 7.470 2.125 ;
        RECT 8.110 2.085 8.280 2.375 ;
        RECT 8.460 2.255 8.840 2.635 ;
        RECT 8.110 1.915 8.960 2.085 ;
        RECT 5.915 1.495 6.690 1.655 ;
        RECT 7.250 1.575 8.620 1.745 ;
        RECT 5.915 0.705 6.125 1.495 ;
        RECT 7.250 1.485 7.470 1.575 ;
        RECT 6.295 0.705 6.745 1.325 ;
        RECT 6.965 1.315 7.470 1.485 ;
        RECT 6.965 0.535 7.135 1.315 ;
        RECT 7.355 0.865 7.625 1.145 ;
        RECT 7.805 1.035 8.395 1.405 ;
        RECT 8.790 1.295 8.960 1.915 ;
        RECT 9.135 1.575 9.305 2.635 ;
        RECT 10.075 1.795 10.245 2.635 ;
        RECT 11.015 1.795 11.185 2.635 ;
        RECT 7.355 0.695 7.935 0.865 ;
        RECT 5.365 0.275 5.765 0.445 ;
        RECT 6.035 0.255 7.135 0.535 ;
        RECT 7.355 0.085 7.595 0.525 ;
        RECT 7.765 0.465 7.935 0.695 ;
        RECT 8.155 0.635 8.395 1.035 ;
        RECT 8.615 1.285 8.960 1.295 ;
        RECT 8.615 1.075 10.795 1.285 ;
        RECT 8.615 0.820 8.940 1.075 ;
        RECT 8.615 0.465 8.935 0.820 ;
        RECT 7.765 0.295 8.935 0.465 ;
        RECT 9.135 0.085 9.305 0.895 ;
        RECT 10.075 0.085 10.245 0.555 ;
        RECT 11.015 0.085 11.185 0.555 ;
        RECT 0.000 -0.085 11.500 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 0.660 1.105 0.830 1.275 ;
        RECT 1.115 1.785 1.285 1.955 ;
        RECT 3.105 1.785 3.275 1.955 ;
        RECT 2.595 1.105 2.765 1.275 ;
        RECT 6.525 1.785 6.695 1.955 ;
        RECT 4.285 0.765 4.455 0.935 ;
        RECT 4.645 0.765 4.815 0.935 ;
        RECT 6.525 1.105 6.695 1.275 ;
        RECT 7.870 1.080 8.040 1.250 ;
        RECT 8.165 0.765 8.335 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
      LAYER met1 ;
        RECT 1.005 1.940 1.345 1.985 ;
        RECT 3.045 1.940 3.335 1.985 ;
        RECT 6.465 1.940 6.805 1.985 ;
        RECT 1.005 1.800 6.805 1.940 ;
        RECT 1.005 1.755 1.345 1.800 ;
        RECT 3.045 1.755 3.335 1.800 ;
        RECT 6.465 1.755 6.805 1.800 ;
        RECT 0.600 1.260 0.890 1.305 ;
        RECT 2.535 1.260 2.825 1.305 ;
        RECT 6.465 1.260 6.805 1.305 ;
        RECT 0.600 1.120 6.805 1.260 ;
        RECT 0.600 1.075 0.890 1.120 ;
        RECT 2.535 1.075 2.825 1.120 ;
        RECT 6.465 1.075 6.805 1.120 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dfrtp_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__dfstp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__dfstp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.120 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.975 0.440 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247200 ;
    PORT
      LAYER li1 ;
        RECT 1.870 1.005 2.330 1.625 ;
    END
  END D
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277200 ;
    PORT
      LAYER met1 ;
        RECT 4.220 0.920 4.510 0.965 ;
        RECT 7.445 0.920 7.735 0.965 ;
        RECT 4.220 0.780 7.735 0.920 ;
        RECT 4.220 0.735 4.510 0.780 ;
        RECT 7.445 0.735 7.735 0.780 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.120 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.465 0.785 2.435 1.005 ;
        RECT 9.095 0.905 10.115 1.015 ;
        RECT 7.580 0.785 10.115 0.905 ;
        RECT 0.005 0.105 10.115 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.310 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.120 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.518250 ;
    PORT
      LAYER li1 ;
        RECT 9.740 1.655 10.025 2.325 ;
        RECT 9.800 0.795 10.025 1.655 ;
        RECT 9.755 0.265 10.025 0.795 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.120 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.895 2.635 ;
        RECT 0.175 1.795 0.890 1.965 ;
        RECT 0.660 0.805 0.890 1.795 ;
        RECT 0.175 0.635 0.890 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.115 0.345 1.340 2.465 ;
        RECT 1.555 2.135 1.885 2.635 ;
        RECT 2.105 1.965 2.275 2.465 ;
        RECT 2.510 2.250 3.440 2.420 ;
        RECT 3.730 2.255 4.110 2.635 ;
        RECT 1.530 1.795 2.275 1.965 ;
        RECT 1.530 0.825 1.700 1.795 ;
        RECT 2.500 1.575 3.100 1.955 ;
        RECT 1.530 0.635 2.275 0.825 ;
        RECT 2.500 0.705 2.770 1.575 ;
        RECT 3.270 1.405 3.440 2.250 ;
        RECT 4.340 2.085 4.510 2.375 ;
        RECT 4.680 2.255 5.060 2.635 ;
        RECT 5.560 2.165 6.290 2.415 ;
        RECT 6.470 2.255 6.940 2.635 ;
        RECT 6.070 2.085 6.290 2.165 ;
        RECT 7.140 2.085 7.380 2.375 ;
        RECT 3.610 1.835 5.110 2.085 ;
        RECT 3.610 1.575 3.910 1.835 ;
        RECT 4.470 1.405 4.770 1.565 ;
        RECT 3.270 1.235 4.770 1.405 ;
        RECT 3.270 1.230 3.740 1.235 ;
        RECT 2.950 0.645 3.350 1.015 ;
        RECT 1.555 0.085 1.885 0.465 ;
        RECT 2.105 0.305 2.275 0.635 ;
        RECT 3.520 0.465 3.740 1.230 ;
        RECT 4.940 1.065 5.110 1.835 ;
        RECT 3.910 0.735 4.510 1.065 ;
        RECT 4.790 0.725 5.110 1.065 ;
        RECT 5.330 1.655 5.900 1.965 ;
        RECT 6.070 1.915 7.380 2.085 ;
        RECT 7.710 1.945 8.040 2.635 ;
        RECT 5.330 0.895 5.500 1.655 ;
        RECT 5.720 1.065 5.900 1.475 ;
        RECT 6.070 1.405 6.290 1.915 ;
        RECT 8.210 1.765 8.380 2.375 ;
        RECT 8.650 1.915 8.980 2.425 ;
        RECT 8.210 1.745 8.550 1.765 ;
        RECT 6.460 1.575 8.550 1.745 ;
        RECT 6.070 1.235 8.170 1.405 ;
        RECT 6.370 0.895 6.750 1.015 ;
        RECT 5.330 0.725 6.750 0.895 ;
        RECT 2.625 0.265 3.740 0.465 ;
        RECT 3.910 0.085 4.370 0.525 ;
        RECT 4.790 0.295 4.960 0.725 ;
        RECT 5.140 0.085 5.530 0.545 ;
        RECT 6.920 0.475 7.090 1.235 ;
        RECT 7.790 1.175 8.170 1.235 ;
        RECT 7.260 1.005 7.640 1.065 ;
        RECT 7.260 0.735 7.780 1.005 ;
        RECT 8.340 0.680 8.550 1.575 ;
        RECT 6.190 0.305 7.090 0.475 ;
        RECT 7.320 0.085 8.030 0.565 ;
        RECT 8.210 0.350 8.550 0.680 ;
        RECT 8.730 1.325 8.980 1.915 ;
        RECT 9.150 1.835 9.570 2.635 ;
        RECT 8.730 0.995 9.580 1.325 ;
        RECT 8.730 0.345 8.980 0.995 ;
        RECT 9.150 0.085 9.585 0.545 ;
        RECT 0.000 -0.085 10.120 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 0.665 1.740 0.835 1.910 ;
        RECT 1.165 0.720 1.335 0.890 ;
        RECT 2.645 1.740 2.815 1.910 ;
        RECT 3.155 0.720 3.325 0.890 ;
        RECT 4.280 0.765 4.450 0.935 ;
        RECT 5.705 1.740 5.875 1.910 ;
        RECT 5.725 1.110 5.895 1.280 ;
        RECT 7.505 0.765 7.675 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
      LAYER met1 ;
        RECT 0.605 1.800 5.935 1.940 ;
        RECT 0.605 1.710 0.895 1.800 ;
        RECT 2.585 1.710 2.875 1.800 ;
        RECT 5.645 1.710 5.935 1.800 ;
        RECT 5.665 1.260 5.955 1.310 ;
        RECT 3.170 1.120 5.955 1.260 ;
        RECT 3.170 0.920 3.385 1.120 ;
        RECT 5.665 1.080 5.955 1.120 ;
        RECT 1.105 0.780 3.385 0.920 ;
        RECT 1.105 0.690 1.395 0.780 ;
        RECT 3.095 0.690 3.385 0.780 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dfstp_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__dfstp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__dfstp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.580 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.975 0.440 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247200 ;
    PORT
      LAYER li1 ;
        RECT 1.870 1.005 2.330 1.625 ;
    END
  END D
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277200 ;
    PORT
      LAYER met1 ;
        RECT 4.220 0.920 4.510 0.965 ;
        RECT 7.445 0.920 7.735 0.965 ;
        RECT 4.220 0.780 7.735 0.920 ;
        RECT 4.220 0.735 4.510 0.780 ;
        RECT 7.445 0.735 7.735 0.780 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.580 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.465 0.785 2.435 1.005 ;
        RECT 8.560 0.905 10.525 1.015 ;
        RECT 7.580 0.785 10.525 0.905 ;
        RECT 0.005 0.105 10.525 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.770 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.580 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.530500 ;
    PORT
      LAYER li1 ;
        RECT 9.540 1.615 10.015 2.460 ;
        RECT 9.540 1.495 10.485 1.615 ;
        RECT 9.750 0.825 10.485 1.495 ;
        RECT 9.685 0.745 10.485 0.825 ;
        RECT 9.685 0.265 10.015 0.745 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.580 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.895 2.635 ;
        RECT 0.175 1.795 0.890 1.965 ;
        RECT 0.660 0.805 0.890 1.795 ;
        RECT 0.175 0.635 0.890 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.115 0.345 1.340 2.465 ;
        RECT 1.555 2.135 1.885 2.635 ;
        RECT 2.105 1.965 2.275 2.465 ;
        RECT 2.510 2.250 3.440 2.420 ;
        RECT 3.730 2.255 4.110 2.635 ;
        RECT 1.530 1.795 2.275 1.965 ;
        RECT 1.530 0.825 1.700 1.795 ;
        RECT 2.500 1.575 3.100 1.955 ;
        RECT 1.530 0.635 2.275 0.825 ;
        RECT 2.500 0.705 2.770 1.575 ;
        RECT 3.270 1.405 3.440 2.250 ;
        RECT 4.340 2.085 4.510 2.375 ;
        RECT 4.680 2.255 5.060 2.635 ;
        RECT 5.560 2.165 6.290 2.415 ;
        RECT 6.470 2.255 6.940 2.635 ;
        RECT 6.070 2.085 6.290 2.165 ;
        RECT 7.140 2.085 7.380 2.375 ;
        RECT 3.610 1.835 5.110 2.085 ;
        RECT 3.610 1.575 3.910 1.835 ;
        RECT 4.470 1.405 4.770 1.565 ;
        RECT 3.270 1.235 4.770 1.405 ;
        RECT 3.270 1.230 3.740 1.235 ;
        RECT 2.950 0.645 3.350 1.015 ;
        RECT 1.555 0.085 1.885 0.465 ;
        RECT 2.105 0.305 2.275 0.635 ;
        RECT 3.520 0.465 3.740 1.230 ;
        RECT 4.940 1.065 5.110 1.835 ;
        RECT 3.910 0.735 4.510 1.065 ;
        RECT 4.790 0.725 5.110 1.065 ;
        RECT 5.330 1.655 5.900 1.965 ;
        RECT 6.070 1.915 7.380 2.085 ;
        RECT 7.710 1.945 8.040 2.635 ;
        RECT 5.330 0.895 5.500 1.655 ;
        RECT 5.720 1.065 5.900 1.475 ;
        RECT 6.070 1.405 6.290 1.915 ;
        RECT 8.210 1.765 8.380 2.375 ;
        RECT 8.650 1.915 8.980 2.425 ;
        RECT 8.210 1.745 8.550 1.765 ;
        RECT 6.460 1.575 8.550 1.745 ;
        RECT 6.070 1.235 8.170 1.405 ;
        RECT 6.370 0.895 6.750 1.015 ;
        RECT 5.330 0.725 6.750 0.895 ;
        RECT 2.625 0.265 3.740 0.465 ;
        RECT 3.910 0.085 4.370 0.525 ;
        RECT 4.790 0.295 4.960 0.725 ;
        RECT 5.140 0.085 5.530 0.545 ;
        RECT 6.920 0.475 7.090 1.235 ;
        RECT 7.790 1.175 8.170 1.235 ;
        RECT 7.260 1.005 7.640 1.065 ;
        RECT 7.260 0.735 7.780 1.005 ;
        RECT 8.340 0.680 8.550 1.575 ;
        RECT 6.190 0.305 7.090 0.475 ;
        RECT 7.320 0.085 8.030 0.565 ;
        RECT 8.210 0.350 8.550 0.680 ;
        RECT 8.730 1.325 8.980 1.915 ;
        RECT 9.200 1.495 9.370 2.635 ;
        RECT 10.185 1.785 10.450 2.635 ;
        RECT 8.730 0.995 9.580 1.325 ;
        RECT 8.730 0.345 8.900 0.995 ;
        RECT 9.070 0.085 9.450 0.825 ;
        RECT 10.185 0.085 10.450 0.575 ;
        RECT 0.000 -0.085 10.580 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 0.665 1.740 0.835 1.910 ;
        RECT 1.165 0.720 1.335 0.890 ;
        RECT 2.645 1.740 2.815 1.910 ;
        RECT 3.155 0.720 3.325 0.890 ;
        RECT 4.280 0.765 4.450 0.935 ;
        RECT 5.705 1.740 5.875 1.910 ;
        RECT 5.725 1.110 5.895 1.280 ;
        RECT 7.505 0.765 7.675 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
      LAYER met1 ;
        RECT 0.605 1.800 5.935 1.940 ;
        RECT 0.605 1.710 0.895 1.800 ;
        RECT 2.585 1.710 2.875 1.800 ;
        RECT 5.645 1.710 5.935 1.800 ;
        RECT 5.665 1.260 5.955 1.310 ;
        RECT 3.170 1.120 5.955 1.260 ;
        RECT 3.170 0.920 3.385 1.120 ;
        RECT 5.665 1.080 5.955 1.120 ;
        RECT 1.105 0.780 3.385 0.920 ;
        RECT 1.105 0.690 1.395 0.780 ;
        RECT 3.095 0.690 3.385 0.780 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dfstp_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__dfstp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__dfstp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.960 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.975 0.440 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247200 ;
    PORT
      LAYER li1 ;
        RECT 1.870 1.005 2.330 1.625 ;
    END
  END D
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277200 ;
    PORT
      LAYER met1 ;
        RECT 4.220 0.920 4.510 0.965 ;
        RECT 7.445 0.920 7.735 0.965 ;
        RECT 4.220 0.780 7.735 0.920 ;
        RECT 4.220 0.735 4.510 0.780 ;
        RECT 7.445 0.735 7.735 0.780 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.960 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.465 0.785 2.435 1.005 ;
        RECT 9.095 0.905 11.945 1.015 ;
        RECT 7.580 0.785 11.945 0.905 ;
        RECT 0.005 0.105 11.945 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 12.150 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.960 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.435000 ;
    PORT
      LAYER li1 ;
        RECT 9.725 1.640 9.995 2.465 ;
        RECT 10.665 1.640 10.835 2.465 ;
        RECT 11.605 1.640 11.860 2.465 ;
        RECT 9.725 1.470 11.860 1.640 ;
        RECT 11.610 0.885 11.860 1.470 ;
        RECT 9.725 0.715 11.860 0.885 ;
        RECT 9.725 0.265 10.025 0.715 ;
        RECT 10.665 0.265 10.835 0.715 ;
        RECT 11.605 0.265 11.860 0.715 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 11.960 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.895 2.635 ;
        RECT 0.175 1.795 0.890 1.965 ;
        RECT 0.660 0.805 0.890 1.795 ;
        RECT 0.175 0.635 0.890 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.115 0.345 1.340 2.465 ;
        RECT 1.555 2.135 1.885 2.635 ;
        RECT 2.105 1.965 2.275 2.465 ;
        RECT 2.510 2.250 3.440 2.420 ;
        RECT 3.730 2.255 4.110 2.635 ;
        RECT 1.530 1.795 2.275 1.965 ;
        RECT 1.530 0.825 1.700 1.795 ;
        RECT 2.500 1.575 3.100 1.955 ;
        RECT 1.530 0.635 2.275 0.825 ;
        RECT 2.500 0.705 2.770 1.575 ;
        RECT 3.270 1.405 3.440 2.250 ;
        RECT 4.340 2.085 4.510 2.375 ;
        RECT 4.680 2.255 5.060 2.635 ;
        RECT 5.560 2.165 6.290 2.415 ;
        RECT 6.470 2.255 6.940 2.635 ;
        RECT 6.070 2.085 6.290 2.165 ;
        RECT 7.140 2.085 7.380 2.375 ;
        RECT 3.610 1.835 5.110 2.085 ;
        RECT 3.610 1.575 3.910 1.835 ;
        RECT 4.470 1.405 4.770 1.565 ;
        RECT 3.270 1.235 4.770 1.405 ;
        RECT 3.270 1.230 3.740 1.235 ;
        RECT 2.950 0.645 3.350 1.015 ;
        RECT 1.555 0.085 1.885 0.465 ;
        RECT 2.105 0.305 2.275 0.635 ;
        RECT 3.520 0.465 3.740 1.230 ;
        RECT 4.940 1.065 5.110 1.835 ;
        RECT 3.910 0.735 4.510 1.065 ;
        RECT 4.790 0.725 5.110 1.065 ;
        RECT 5.330 1.655 5.900 1.965 ;
        RECT 6.070 1.915 7.380 2.085 ;
        RECT 7.710 1.945 8.040 2.635 ;
        RECT 5.330 0.895 5.500 1.655 ;
        RECT 5.720 1.065 5.900 1.475 ;
        RECT 6.070 1.405 6.290 1.915 ;
        RECT 8.210 1.765 8.380 2.375 ;
        RECT 8.650 1.915 8.980 2.425 ;
        RECT 8.210 1.745 8.550 1.765 ;
        RECT 6.460 1.575 8.550 1.745 ;
        RECT 6.070 1.235 8.170 1.405 ;
        RECT 6.370 0.895 6.750 1.015 ;
        RECT 5.330 0.725 6.750 0.895 ;
        RECT 2.625 0.265 3.740 0.465 ;
        RECT 3.910 0.085 4.370 0.525 ;
        RECT 4.790 0.295 4.960 0.725 ;
        RECT 5.140 0.085 5.530 0.545 ;
        RECT 6.920 0.475 7.090 1.235 ;
        RECT 7.790 1.175 8.170 1.235 ;
        RECT 7.260 1.005 7.640 1.065 ;
        RECT 7.260 0.735 7.780 1.005 ;
        RECT 8.340 0.680 8.550 1.575 ;
        RECT 6.190 0.305 7.090 0.475 ;
        RECT 7.320 0.085 8.030 0.565 ;
        RECT 8.210 0.350 8.550 0.680 ;
        RECT 8.730 1.275 8.980 1.915 ;
        RECT 9.190 1.835 9.545 2.635 ;
        RECT 10.165 1.810 10.420 2.635 ;
        RECT 11.055 1.810 11.435 2.635 ;
        RECT 8.730 1.055 11.440 1.275 ;
        RECT 8.730 0.345 8.980 1.055 ;
        RECT 9.190 0.085 9.475 0.545 ;
        RECT 10.195 0.085 10.495 0.545 ;
        RECT 11.055 0.085 11.435 0.545 ;
        RECT 0.000 -0.085 11.960 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 0.665 1.740 0.835 1.910 ;
        RECT 1.165 0.720 1.335 0.890 ;
        RECT 2.645 1.740 2.815 1.910 ;
        RECT 3.155 0.720 3.325 0.890 ;
        RECT 4.280 0.765 4.450 0.935 ;
        RECT 5.705 1.740 5.875 1.910 ;
        RECT 5.725 1.110 5.895 1.280 ;
        RECT 7.505 0.765 7.675 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
      LAYER met1 ;
        RECT 0.605 1.800 5.935 1.940 ;
        RECT 0.605 1.710 0.895 1.800 ;
        RECT 2.585 1.710 2.875 1.800 ;
        RECT 5.645 1.710 5.935 1.800 ;
        RECT 5.665 1.260 5.955 1.310 ;
        RECT 3.170 1.120 5.955 1.260 ;
        RECT 3.170 0.920 3.385 1.120 ;
        RECT 5.665 1.080 5.955 1.120 ;
        RECT 1.105 0.780 3.385 0.920 ;
        RECT 1.105 0.690 1.395 0.780 ;
        RECT 3.095 0.690 3.385 0.780 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dfstp_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__diode_2
  CLASS CORE ANTENNACELL ;
  FOREIGN sky130_fd_sc_hdll__diode_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.920 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN DIODE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.835 2.465 ;
    END
  END DIODE
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 0.920 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.025 0.065 0.915 1.015 ;
        RECT 0.145 -0.085 0.315 0.065 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 1.110 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 0.920 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 0.920 2.805 ;
        RECT 0.000 -0.085 0.920 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__diode_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__diode_4
  CLASS CORE ANTENNACELL ;
  FOREIGN sky130_fd_sc_hdll__diode_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN DIODE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.055700 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 1.755 2.465 ;
    END
  END DIODE
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.025 0.065 1.815 1.015 ;
        RECT 0.145 -0.085 0.315 0.065 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.840 2.805 ;
        RECT 0.000 -0.085 1.840 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__diode_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__diode_6
  CLASS CORE ANTENNACELL ;
  FOREIGN sky130_fd_sc_hdll__diode_6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN DIODE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.203200 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 2.675 2.465 ;
    END
  END DIODE
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.935 1.015 1.825 1.785 ;
        RECT 0.005 0.065 2.755 1.015 ;
        RECT 0.145 -0.085 0.315 0.065 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 2.070 2.950 2.910 ;
        RECT -0.190 1.305 0.650 2.070 ;
        RECT 2.110 1.305 2.950 2.070 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__diode_6

#--------EOF---------

MACRO sky130_fd_sc_hdll__diode_8
  CLASS CORE ANTENNACELL ;
  FOREIGN sky130_fd_sc_hdll__diode_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN DIODE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.546400 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 3.595 2.465 ;
    END
  END DIODE
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.935 1.015 2.745 1.785 ;
        RECT 0.005 0.065 3.675 1.015 ;
        RECT 0.145 -0.085 0.315 0.065 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 2.070 3.870 2.910 ;
        RECT -0.190 1.305 0.650 2.070 ;
        RECT 3.030 1.305 3.870 2.070 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__diode_8

#--------EOF---------

MACRO sky130_fd_sc_hdll__dlrtn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__dlrtn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 1.435 0.955 1.765 1.300 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.435 1.625 ;
    END
  END GATE_N
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 4.890 0.995 5.385 1.325 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.365 0.785 6.185 1.015 ;
        RECT 0.055 0.105 6.185 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 5.815 2.255 6.295 2.465 ;
        RECT 5.895 1.495 6.295 2.255 ;
        RECT 6.065 0.885 6.295 1.495 ;
        RECT 5.820 0.495 6.295 0.885 ;
        RECT 5.765 0.255 6.295 0.495 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.085 1.965 0.395 2.465 ;
        RECT 0.565 2.135 0.895 2.635 ;
        RECT 0.085 1.795 0.895 1.965 ;
        RECT 0.605 1.070 0.895 1.795 ;
        RECT 1.065 1.445 1.335 2.465 ;
        RECT 1.555 1.665 1.885 2.465 ;
        RECT 2.055 1.835 2.325 2.635 ;
        RECT 3.020 2.165 3.850 2.385 ;
        RECT 1.555 1.495 2.115 1.665 ;
        RECT 0.605 0.805 0.775 1.070 ;
        RECT 0.225 0.635 0.775 0.805 ;
        RECT 0.225 0.280 0.395 0.635 ;
        RECT 0.565 0.085 0.895 0.465 ;
        RECT 1.065 0.280 1.235 1.445 ;
        RECT 1.945 1.095 2.115 1.495 ;
        RECT 2.445 1.265 2.955 1.685 ;
        RECT 3.125 1.575 3.510 1.995 ;
        RECT 3.125 1.095 3.295 1.575 ;
        RECT 3.680 1.325 3.850 2.165 ;
        RECT 4.050 2.135 4.635 2.635 ;
        RECT 4.885 1.865 5.170 2.465 ;
        RECT 5.345 2.150 5.645 2.635 ;
        RECT 5.345 1.885 5.675 2.150 ;
        RECT 4.020 1.705 5.170 1.865 ;
        RECT 4.020 1.535 5.725 1.705 ;
        RECT 3.680 1.165 4.380 1.325 ;
        RECT 1.945 0.785 2.535 1.095 ;
        RECT 1.660 0.765 2.535 0.785 ;
        RECT 1.660 0.615 2.115 0.765 ;
        RECT 2.780 0.735 3.295 1.095 ;
        RECT 3.490 0.995 4.380 1.165 ;
        RECT 1.660 0.345 1.855 0.615 ;
        RECT 3.490 0.565 3.660 0.995 ;
        RECT 4.550 0.825 4.720 1.535 ;
        RECT 5.555 1.325 5.725 1.535 ;
        RECT 5.555 1.055 5.895 1.325 ;
        RECT 2.025 0.085 2.355 0.445 ;
        RECT 3.040 0.280 3.660 0.565 ;
        RECT 3.870 0.085 4.200 0.610 ;
        RECT 4.455 0.255 4.785 0.825 ;
        RECT 5.320 0.625 5.650 0.825 ;
        RECT 5.320 0.085 5.595 0.625 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.635 1.785 0.805 1.955 ;
        RECT 1.095 1.445 1.265 1.615 ;
        RECT 3.280 1.785 3.450 1.955 ;
        RECT 2.725 1.445 2.895 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
      LAYER met1 ;
        RECT 0.575 1.940 0.865 1.985 ;
        RECT 3.220 1.940 3.510 1.985 ;
        RECT 0.575 1.800 3.510 1.940 ;
        RECT 0.575 1.755 0.865 1.800 ;
        RECT 3.220 1.755 3.510 1.800 ;
        RECT 1.035 1.600 1.325 1.645 ;
        RECT 2.665 1.600 2.955 1.645 ;
        RECT 1.035 1.460 2.955 1.600 ;
        RECT 1.035 1.415 1.325 1.460 ;
        RECT 2.665 1.415 2.955 1.460 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dlrtn_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__dlrtn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__dlrtn_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.900 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 1.435 0.955 1.765 1.300 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.435 1.625 ;
    END
  END GATE_N
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 4.890 0.995 5.385 1.325 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.900 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.365 0.785 6.715 1.015 ;
        RECT 0.055 0.105 6.715 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.090 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.900 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.465500 ;
    PORT
      LAYER li1 ;
        RECT 5.815 2.255 6.205 2.455 ;
        RECT 5.895 1.495 6.205 2.255 ;
        RECT 6.035 1.325 6.205 1.495 ;
        RECT 6.035 1.055 6.435 1.325 ;
        RECT 6.035 0.825 6.205 1.055 ;
        RECT 5.815 0.255 6.205 0.825 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.900 2.805 ;
        RECT 0.085 1.965 0.395 2.465 ;
        RECT 0.565 2.135 0.895 2.635 ;
        RECT 0.085 1.795 0.895 1.965 ;
        RECT 0.605 1.070 0.895 1.795 ;
        RECT 1.065 1.445 1.335 2.465 ;
        RECT 1.555 1.665 1.885 2.465 ;
        RECT 2.055 1.835 2.325 2.635 ;
        RECT 3.020 2.165 3.850 2.385 ;
        RECT 1.555 1.495 2.115 1.665 ;
        RECT 0.605 0.805 0.775 1.070 ;
        RECT 0.225 0.635 0.775 0.805 ;
        RECT 0.225 0.280 0.395 0.635 ;
        RECT 0.565 0.085 0.895 0.465 ;
        RECT 1.065 0.280 1.235 1.445 ;
        RECT 1.945 1.095 2.115 1.495 ;
        RECT 2.445 1.265 2.955 1.685 ;
        RECT 3.125 1.575 3.510 1.995 ;
        RECT 3.125 1.095 3.295 1.575 ;
        RECT 3.680 1.325 3.850 2.165 ;
        RECT 4.050 2.135 4.635 2.635 ;
        RECT 4.885 1.865 5.170 2.465 ;
        RECT 5.345 2.150 5.645 2.635 ;
        RECT 5.345 1.885 5.675 2.150 ;
        RECT 4.020 1.705 5.170 1.865 ;
        RECT 4.020 1.535 5.725 1.705 ;
        RECT 3.680 1.165 4.380 1.325 ;
        RECT 1.945 0.785 2.535 1.095 ;
        RECT 1.660 0.765 2.535 0.785 ;
        RECT 1.660 0.615 2.115 0.765 ;
        RECT 2.780 0.735 3.295 1.095 ;
        RECT 3.490 0.995 4.380 1.165 ;
        RECT 1.660 0.345 1.855 0.615 ;
        RECT 3.490 0.565 3.660 0.995 ;
        RECT 4.550 0.825 4.720 1.535 ;
        RECT 5.555 1.325 5.725 1.535 ;
        RECT 6.375 1.495 6.580 2.635 ;
        RECT 5.555 0.995 5.865 1.325 ;
        RECT 2.025 0.085 2.355 0.445 ;
        RECT 3.040 0.280 3.660 0.565 ;
        RECT 3.870 0.085 4.200 0.610 ;
        RECT 4.455 0.255 4.785 0.825 ;
        RECT 5.315 0.085 5.645 0.825 ;
        RECT 6.375 0.085 6.585 0.885 ;
        RECT 0.000 -0.085 6.900 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 0.635 1.785 0.805 1.955 ;
        RECT 1.095 1.445 1.265 1.615 ;
        RECT 3.280 1.785 3.450 1.955 ;
        RECT 2.725 1.445 2.895 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
      LAYER met1 ;
        RECT 0.575 1.940 0.865 1.985 ;
        RECT 3.220 1.940 3.510 1.985 ;
        RECT 0.575 1.800 3.510 1.940 ;
        RECT 0.575 1.755 0.865 1.800 ;
        RECT 3.220 1.755 3.510 1.800 ;
        RECT 1.035 1.600 1.325 1.645 ;
        RECT 2.665 1.600 2.955 1.645 ;
        RECT 1.035 1.460 2.955 1.600 ;
        RECT 1.035 1.415 1.325 1.460 ;
        RECT 2.665 1.415 2.955 1.460 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dlrtn_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__dlrtn_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__dlrtn_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.820 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 1.435 0.955 1.765 1.300 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.435 1.625 ;
    END
  END GATE_N
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 4.890 0.995 5.385 1.325 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.820 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.365 0.785 7.595 1.015 ;
        RECT 0.055 0.105 7.595 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.010 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.820 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.931000 ;
    PORT
      LAYER li1 ;
        RECT 5.815 2.255 6.145 2.465 ;
        RECT 5.845 1.875 6.145 2.255 ;
        RECT 5.895 1.665 6.145 1.875 ;
        RECT 6.755 1.665 7.085 2.465 ;
        RECT 5.895 1.495 7.085 1.665 ;
        RECT 6.405 1.325 7.085 1.495 ;
        RECT 6.405 1.055 7.265 1.325 ;
        RECT 6.405 0.905 7.085 1.055 ;
        RECT 5.815 0.735 7.085 0.905 ;
        RECT 5.815 0.255 6.195 0.735 ;
        RECT 6.755 0.255 7.085 0.735 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.820 2.805 ;
        RECT 0.085 1.965 0.395 2.465 ;
        RECT 0.565 2.135 0.895 2.635 ;
        RECT 0.085 1.795 0.895 1.965 ;
        RECT 0.605 1.070 0.895 1.795 ;
        RECT 1.065 1.445 1.335 2.465 ;
        RECT 1.555 1.665 1.885 2.465 ;
        RECT 2.055 1.835 2.325 2.635 ;
        RECT 3.020 2.165 3.850 2.385 ;
        RECT 1.555 1.495 2.115 1.665 ;
        RECT 0.605 0.805 0.775 1.070 ;
        RECT 0.225 0.635 0.775 0.805 ;
        RECT 0.225 0.280 0.395 0.635 ;
        RECT 0.565 0.085 0.895 0.465 ;
        RECT 1.065 0.280 1.235 1.445 ;
        RECT 1.945 1.095 2.115 1.495 ;
        RECT 2.445 1.265 2.955 1.685 ;
        RECT 3.125 1.575 3.510 1.995 ;
        RECT 3.125 1.095 3.295 1.575 ;
        RECT 3.680 1.325 3.850 2.165 ;
        RECT 4.020 2.135 4.705 2.635 ;
        RECT 4.875 1.865 5.175 2.435 ;
        RECT 5.345 2.150 5.645 2.635 ;
        RECT 5.345 1.875 5.675 2.150 ;
        RECT 4.020 1.705 5.175 1.865 ;
        RECT 6.315 1.835 6.585 2.635 ;
        RECT 4.020 1.535 5.725 1.705 ;
        RECT 3.680 1.165 4.380 1.325 ;
        RECT 1.945 0.785 2.535 1.095 ;
        RECT 1.660 0.765 2.535 0.785 ;
        RECT 1.660 0.615 2.115 0.765 ;
        RECT 2.780 0.735 3.295 1.095 ;
        RECT 3.490 0.995 4.380 1.165 ;
        RECT 1.660 0.345 1.855 0.615 ;
        RECT 3.490 0.565 3.660 0.995 ;
        RECT 4.550 0.825 4.720 1.535 ;
        RECT 5.555 1.325 5.725 1.535 ;
        RECT 7.255 1.495 7.510 2.635 ;
        RECT 5.555 1.075 6.235 1.325 ;
        RECT 2.025 0.085 2.355 0.445 ;
        RECT 3.040 0.280 3.660 0.565 ;
        RECT 3.870 0.085 4.200 0.610 ;
        RECT 4.455 0.255 4.785 0.825 ;
        RECT 5.315 0.085 5.645 0.825 ;
        RECT 6.375 0.085 6.585 0.565 ;
        RECT 7.255 0.085 7.465 0.885 ;
        RECT 0.000 -0.085 7.820 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 0.635 1.785 0.805 1.955 ;
        RECT 1.095 1.445 1.265 1.615 ;
        RECT 3.280 1.785 3.450 1.955 ;
        RECT 2.725 1.445 2.895 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
      LAYER met1 ;
        RECT 0.575 1.940 0.865 1.985 ;
        RECT 3.220 1.940 3.510 1.985 ;
        RECT 0.575 1.800 3.510 1.940 ;
        RECT 0.575 1.755 0.865 1.800 ;
        RECT 3.220 1.755 3.510 1.800 ;
        RECT 1.035 1.600 1.325 1.645 ;
        RECT 2.665 1.600 2.955 1.645 ;
        RECT 1.035 1.460 2.955 1.600 ;
        RECT 1.035 1.415 1.325 1.460 ;
        RECT 2.665 1.415 2.955 1.460 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dlrtn_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__dlrtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__dlrtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 1.435 0.955 1.765 1.325 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.435 1.625 ;
    END
  END GATE
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 4.890 0.995 5.385 1.325 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.365 0.785 6.185 1.015 ;
        RECT 0.055 0.105 6.185 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 5.815 2.255 6.295 2.465 ;
        RECT 5.895 1.495 6.295 2.255 ;
        RECT 6.065 0.885 6.295 1.495 ;
        RECT 5.820 0.495 6.295 0.885 ;
        RECT 5.765 0.255 6.295 0.495 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.085 1.965 0.395 2.465 ;
        RECT 0.565 2.135 0.895 2.635 ;
        RECT 0.085 1.795 0.775 1.965 ;
        RECT 0.605 1.400 0.775 1.795 ;
        RECT 1.065 1.685 1.335 2.465 ;
        RECT 0.605 1.070 0.895 1.400 ;
        RECT 0.605 0.805 0.775 1.070 ;
        RECT 0.225 0.635 0.775 0.805 ;
        RECT 0.225 0.280 0.395 0.635 ;
        RECT 0.565 0.085 0.895 0.465 ;
        RECT 1.065 0.280 1.235 1.685 ;
        RECT 1.555 1.665 1.885 2.465 ;
        RECT 2.055 1.835 2.325 2.635 ;
        RECT 3.020 2.165 3.850 2.385 ;
        RECT 1.555 1.495 2.115 1.665 ;
        RECT 1.945 1.095 2.115 1.495 ;
        RECT 2.445 1.265 2.955 1.685 ;
        RECT 3.125 1.575 3.510 1.995 ;
        RECT 3.125 1.095 3.295 1.575 ;
        RECT 3.680 1.325 3.850 2.165 ;
        RECT 4.050 2.135 4.635 2.635 ;
        RECT 4.885 1.865 5.170 2.465 ;
        RECT 5.345 2.150 5.645 2.635 ;
        RECT 5.345 1.885 5.675 2.150 ;
        RECT 4.020 1.705 5.170 1.865 ;
        RECT 4.020 1.535 5.725 1.705 ;
        RECT 3.680 1.165 4.380 1.325 ;
        RECT 1.945 0.785 2.535 1.095 ;
        RECT 1.660 0.765 2.535 0.785 ;
        RECT 1.660 0.615 2.115 0.765 ;
        RECT 2.780 0.735 3.295 1.095 ;
        RECT 3.490 0.995 4.380 1.165 ;
        RECT 1.660 0.345 1.855 0.615 ;
        RECT 3.490 0.565 3.660 0.995 ;
        RECT 4.550 0.825 4.720 1.535 ;
        RECT 5.555 1.325 5.725 1.535 ;
        RECT 5.555 1.055 5.895 1.325 ;
        RECT 2.025 0.085 2.355 0.445 ;
        RECT 3.040 0.280 3.660 0.565 ;
        RECT 3.870 0.085 4.200 0.610 ;
        RECT 4.455 0.255 4.785 0.825 ;
        RECT 5.320 0.625 5.650 0.825 ;
        RECT 5.320 0.085 5.595 0.625 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.605 1.445 0.775 1.615 ;
        RECT 1.115 1.785 1.285 1.955 ;
        RECT 3.280 1.785 3.450 1.955 ;
        RECT 2.725 1.445 2.895 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
      LAYER met1 ;
        RECT 1.055 1.940 1.345 1.985 ;
        RECT 3.220 1.940 3.510 1.985 ;
        RECT 1.055 1.800 3.510 1.940 ;
        RECT 1.055 1.755 1.345 1.800 ;
        RECT 3.220 1.755 3.510 1.800 ;
        RECT 0.545 1.600 0.835 1.645 ;
        RECT 2.665 1.600 2.955 1.645 ;
        RECT 0.545 1.460 2.955 1.600 ;
        RECT 0.545 1.415 0.835 1.460 ;
        RECT 2.665 1.415 2.955 1.460 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dlrtp_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__dlrtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__dlrtp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.900 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 1.435 0.955 1.765 1.325 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.435 1.625 ;
    END
  END GATE
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 4.890 0.995 5.385 1.325 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.900 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.365 0.785 6.715 1.015 ;
        RECT 0.055 0.105 6.715 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.090 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.900 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.465500 ;
    PORT
      LAYER li1 ;
        RECT 5.815 2.255 6.205 2.455 ;
        RECT 5.895 1.495 6.205 2.255 ;
        RECT 6.035 1.325 6.205 1.495 ;
        RECT 6.035 1.055 6.435 1.325 ;
        RECT 6.035 0.825 6.205 1.055 ;
        RECT 5.815 0.255 6.205 0.825 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.900 2.805 ;
        RECT 0.085 1.965 0.395 2.465 ;
        RECT 0.565 2.135 0.895 2.635 ;
        RECT 0.085 1.795 0.775 1.965 ;
        RECT 0.605 1.400 0.775 1.795 ;
        RECT 1.065 1.685 1.335 2.465 ;
        RECT 0.605 1.070 0.895 1.400 ;
        RECT 0.605 0.805 0.775 1.070 ;
        RECT 0.225 0.635 0.775 0.805 ;
        RECT 0.225 0.280 0.395 0.635 ;
        RECT 0.565 0.085 0.895 0.465 ;
        RECT 1.065 0.280 1.235 1.685 ;
        RECT 1.555 1.665 1.885 2.465 ;
        RECT 2.055 1.835 2.325 2.635 ;
        RECT 3.020 2.165 3.850 2.385 ;
        RECT 1.555 1.495 2.115 1.665 ;
        RECT 1.945 1.095 2.115 1.495 ;
        RECT 2.445 1.265 2.955 1.685 ;
        RECT 3.125 1.575 3.510 1.995 ;
        RECT 3.125 1.095 3.295 1.575 ;
        RECT 3.680 1.325 3.850 2.165 ;
        RECT 4.050 2.135 4.635 2.635 ;
        RECT 4.885 1.865 5.170 2.465 ;
        RECT 5.345 2.150 5.645 2.635 ;
        RECT 5.345 1.885 5.675 2.150 ;
        RECT 4.020 1.705 5.170 1.865 ;
        RECT 4.020 1.535 5.725 1.705 ;
        RECT 3.680 1.165 4.380 1.325 ;
        RECT 1.945 0.785 2.535 1.095 ;
        RECT 1.660 0.765 2.535 0.785 ;
        RECT 1.660 0.615 2.115 0.765 ;
        RECT 2.780 0.735 3.295 1.095 ;
        RECT 3.490 0.995 4.380 1.165 ;
        RECT 1.660 0.345 1.855 0.615 ;
        RECT 3.490 0.565 3.660 0.995 ;
        RECT 4.550 0.825 4.720 1.535 ;
        RECT 5.555 1.325 5.725 1.535 ;
        RECT 6.375 1.495 6.580 2.635 ;
        RECT 5.555 0.995 5.865 1.325 ;
        RECT 2.025 0.085 2.355 0.445 ;
        RECT 3.040 0.280 3.660 0.565 ;
        RECT 3.870 0.085 4.200 0.610 ;
        RECT 4.455 0.255 4.785 0.825 ;
        RECT 5.315 0.085 5.645 0.825 ;
        RECT 6.375 0.085 6.585 0.885 ;
        RECT 0.000 -0.085 6.900 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 0.605 1.445 0.775 1.615 ;
        RECT 1.115 1.785 1.285 1.955 ;
        RECT 3.280 1.785 3.450 1.955 ;
        RECT 2.725 1.445 2.895 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
      LAYER met1 ;
        RECT 1.055 1.940 1.345 1.985 ;
        RECT 3.220 1.940 3.510 1.985 ;
        RECT 1.055 1.800 3.510 1.940 ;
        RECT 1.055 1.755 1.345 1.800 ;
        RECT 3.220 1.755 3.510 1.800 ;
        RECT 0.545 1.600 0.835 1.645 ;
        RECT 2.665 1.600 2.955 1.645 ;
        RECT 0.545 1.460 2.955 1.600 ;
        RECT 0.545 1.415 0.835 1.460 ;
        RECT 2.665 1.415 2.955 1.460 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dlrtp_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__dlrtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__dlrtp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.820 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 1.435 0.955 1.765 1.325 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.435 1.625 ;
    END
  END GATE
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 4.890 0.995 5.385 1.325 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.820 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.365 0.785 7.595 1.015 ;
        RECT 0.055 0.105 7.595 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.010 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.820 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.931000 ;
    PORT
      LAYER li1 ;
        RECT 5.815 2.255 6.145 2.465 ;
        RECT 5.845 1.875 6.145 2.255 ;
        RECT 5.895 1.665 6.145 1.875 ;
        RECT 6.755 1.665 7.085 2.465 ;
        RECT 5.895 1.495 7.085 1.665 ;
        RECT 6.405 1.325 7.085 1.495 ;
        RECT 6.405 1.055 7.265 1.325 ;
        RECT 6.405 0.905 7.085 1.055 ;
        RECT 5.815 0.735 7.085 0.905 ;
        RECT 5.815 0.255 6.195 0.735 ;
        RECT 6.755 0.255 7.085 0.735 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.820 2.805 ;
        RECT 0.085 1.965 0.395 2.465 ;
        RECT 0.565 2.135 0.895 2.635 ;
        RECT 0.085 1.795 0.775 1.965 ;
        RECT 0.605 1.400 0.775 1.795 ;
        RECT 1.065 1.685 1.335 2.465 ;
        RECT 0.605 1.070 0.895 1.400 ;
        RECT 0.605 0.805 0.775 1.070 ;
        RECT 0.225 0.635 0.775 0.805 ;
        RECT 0.225 0.280 0.395 0.635 ;
        RECT 0.565 0.085 0.895 0.465 ;
        RECT 1.065 0.280 1.235 1.685 ;
        RECT 1.555 1.665 1.885 2.465 ;
        RECT 2.055 1.835 2.325 2.635 ;
        RECT 3.020 2.165 3.850 2.385 ;
        RECT 1.555 1.495 2.115 1.665 ;
        RECT 1.945 1.095 2.115 1.495 ;
        RECT 2.445 1.265 2.955 1.685 ;
        RECT 3.125 1.575 3.510 1.995 ;
        RECT 3.125 1.095 3.295 1.575 ;
        RECT 3.680 1.325 3.850 2.165 ;
        RECT 4.020 2.135 4.705 2.635 ;
        RECT 4.875 1.865 5.175 2.435 ;
        RECT 5.345 2.150 5.645 2.635 ;
        RECT 5.345 1.875 5.675 2.150 ;
        RECT 4.020 1.705 5.175 1.865 ;
        RECT 6.315 1.835 6.585 2.635 ;
        RECT 4.020 1.535 5.725 1.705 ;
        RECT 3.680 1.165 4.380 1.325 ;
        RECT 1.945 0.785 2.535 1.095 ;
        RECT 1.660 0.765 2.535 0.785 ;
        RECT 1.660 0.615 2.115 0.765 ;
        RECT 2.780 0.735 3.295 1.095 ;
        RECT 3.490 0.995 4.380 1.165 ;
        RECT 1.660 0.345 1.855 0.615 ;
        RECT 3.490 0.565 3.660 0.995 ;
        RECT 4.550 0.825 4.720 1.535 ;
        RECT 5.555 1.325 5.725 1.535 ;
        RECT 7.255 1.495 7.510 2.635 ;
        RECT 5.555 1.075 6.235 1.325 ;
        RECT 2.025 0.085 2.355 0.445 ;
        RECT 3.040 0.280 3.660 0.565 ;
        RECT 3.870 0.085 4.200 0.610 ;
        RECT 4.455 0.255 4.785 0.825 ;
        RECT 5.315 0.085 5.645 0.825 ;
        RECT 6.375 0.085 6.585 0.565 ;
        RECT 7.255 0.085 7.465 0.885 ;
        RECT 0.000 -0.085 7.820 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 0.605 1.445 0.775 1.615 ;
        RECT 1.115 1.785 1.285 1.955 ;
        RECT 3.280 1.785 3.450 1.955 ;
        RECT 2.725 1.445 2.895 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
      LAYER met1 ;
        RECT 1.055 1.940 1.345 1.985 ;
        RECT 3.220 1.940 3.510 1.985 ;
        RECT 1.055 1.800 3.510 1.940 ;
        RECT 1.055 1.755 1.345 1.800 ;
        RECT 3.220 1.755 3.510 1.800 ;
        RECT 0.545 1.600 0.835 1.645 ;
        RECT 2.665 1.600 2.955 1.645 ;
        RECT 0.545 1.460 2.955 1.600 ;
        RECT 0.545 1.415 0.835 1.460 ;
        RECT 2.665 1.415 2.955 1.460 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dlrtp_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__dlxtn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__dlxtn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 1.465 0.955 1.890 1.325 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.330 1.625 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.400 0.785 5.930 1.015 ;
        RECT 0.005 0.105 5.930 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.554500 ;
    PORT
      LAYER li1 ;
        RECT 5.590 0.415 5.875 2.455 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.895 2.635 ;
        RECT 0.175 1.795 0.830 1.965 ;
        RECT 0.660 1.400 0.830 1.795 ;
        RECT 1.115 1.685 1.340 2.465 ;
        RECT 0.660 1.070 0.890 1.400 ;
        RECT 0.660 0.805 0.830 1.070 ;
        RECT 0.175 0.635 0.830 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.115 0.345 1.285 1.685 ;
        RECT 1.555 1.665 1.885 2.415 ;
        RECT 2.105 1.835 2.420 2.635 ;
        RECT 3.020 2.255 3.850 2.425 ;
        RECT 1.555 1.495 2.290 1.665 ;
        RECT 2.120 1.095 2.290 1.495 ;
        RECT 2.670 1.355 2.955 2.005 ;
        RECT 3.170 1.415 3.510 1.995 ;
        RECT 2.120 0.785 2.540 1.095 ;
        RECT 3.170 1.035 3.340 1.415 ;
        RECT 1.635 0.765 2.540 0.785 ;
        RECT 1.635 0.615 2.290 0.765 ;
        RECT 2.885 0.705 3.340 1.035 ;
        RECT 3.680 1.325 3.850 2.255 ;
        RECT 4.050 2.135 4.350 2.635 ;
        RECT 4.570 1.865 4.790 2.435 ;
        RECT 4.070 1.535 4.790 1.865 ;
        RECT 4.620 1.325 4.790 1.535 ;
        RECT 5.020 1.495 5.290 2.635 ;
        RECT 3.680 0.995 4.430 1.325 ;
        RECT 4.620 0.995 5.420 1.325 ;
        RECT 1.635 0.345 1.805 0.615 ;
        RECT 3.680 0.535 3.850 0.995 ;
        RECT 4.620 0.825 4.790 0.995 ;
        RECT 1.975 0.085 2.355 0.445 ;
        RECT 3.005 0.365 3.850 0.535 ;
        RECT 4.020 0.085 4.300 0.825 ;
        RECT 4.570 0.415 4.790 0.825 ;
        RECT 5.020 0.085 5.290 0.825 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.660 1.445 0.830 1.615 ;
        RECT 1.170 1.785 1.340 1.955 ;
        RECT 2.670 1.785 2.840 1.955 ;
        RECT 3.175 1.445 3.345 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
      LAYER met1 ;
        RECT 1.110 1.940 1.400 1.985 ;
        RECT 2.610 1.940 2.900 1.985 ;
        RECT 1.110 1.800 2.900 1.940 ;
        RECT 1.110 1.755 1.400 1.800 ;
        RECT 2.610 1.755 2.900 1.800 ;
        RECT 0.600 1.600 0.890 1.645 ;
        RECT 3.115 1.600 3.405 1.645 ;
        RECT 0.600 1.460 3.405 1.600 ;
        RECT 0.600 1.415 0.890 1.460 ;
        RECT 3.115 1.415 3.405 1.460 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dlxtn_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__dlxtn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__dlxtn_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 1.465 0.955 1.890 1.325 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.330 1.625 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.515 0.785 6.435 1.015 ;
        RECT 0.005 0.105 6.435 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.498000 ;
    PORT
      LAYER li1 ;
        RECT 5.625 1.495 5.910 2.455 ;
        RECT 5.740 1.325 5.910 1.495 ;
        RECT 5.740 0.995 6.345 1.325 ;
        RECT 5.740 0.825 5.910 0.995 ;
        RECT 5.625 0.415 5.910 0.825 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.895 2.635 ;
        RECT 0.175 1.795 0.830 1.965 ;
        RECT 0.660 1.400 0.830 1.795 ;
        RECT 1.115 1.685 1.340 2.465 ;
        RECT 0.660 1.070 0.890 1.400 ;
        RECT 0.660 0.805 0.830 1.070 ;
        RECT 0.175 0.635 0.830 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.115 0.345 1.285 1.685 ;
        RECT 1.555 1.665 1.885 2.415 ;
        RECT 2.105 1.835 2.420 2.635 ;
        RECT 3.145 2.255 3.945 2.425 ;
        RECT 1.555 1.495 2.290 1.665 ;
        RECT 2.120 1.095 2.290 1.495 ;
        RECT 2.670 1.355 2.955 2.005 ;
        RECT 3.170 1.415 3.510 1.995 ;
        RECT 2.120 0.785 2.540 1.095 ;
        RECT 3.170 1.035 3.340 1.415 ;
        RECT 3.775 1.325 3.945 2.255 ;
        RECT 4.165 2.135 4.465 2.635 ;
        RECT 4.685 1.865 4.905 2.435 ;
        RECT 4.185 1.535 4.905 1.865 ;
        RECT 4.735 1.325 4.905 1.535 ;
        RECT 5.135 1.495 5.405 2.635 ;
        RECT 6.095 1.755 6.345 2.635 ;
        RECT 3.775 1.165 4.545 1.325 ;
        RECT 1.635 0.765 2.540 0.785 ;
        RECT 1.635 0.615 2.290 0.765 ;
        RECT 2.915 0.705 3.340 1.035 ;
        RECT 3.625 0.995 4.545 1.165 ;
        RECT 4.735 0.995 5.535 1.325 ;
        RECT 1.635 0.345 1.805 0.615 ;
        RECT 3.625 0.535 3.795 0.995 ;
        RECT 4.735 0.825 4.905 0.995 ;
        RECT 1.975 0.085 2.355 0.445 ;
        RECT 3.085 0.365 3.795 0.535 ;
        RECT 4.035 0.085 4.415 0.825 ;
        RECT 4.685 0.415 4.905 0.825 ;
        RECT 5.135 0.085 5.405 0.825 ;
        RECT 6.095 0.085 6.355 0.550 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.660 1.445 0.830 1.615 ;
        RECT 1.170 1.785 1.340 1.955 ;
        RECT 2.670 1.785 2.840 1.955 ;
        RECT 3.175 1.445 3.345 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
      LAYER met1 ;
        RECT 1.110 1.940 1.400 1.985 ;
        RECT 2.610 1.940 2.900 1.985 ;
        RECT 1.110 1.800 2.900 1.940 ;
        RECT 1.110 1.755 1.400 1.800 ;
        RECT 2.610 1.755 2.900 1.800 ;
        RECT 0.600 1.600 0.890 1.645 ;
        RECT 3.115 1.600 3.405 1.645 ;
        RECT 0.600 1.460 3.405 1.600 ;
        RECT 0.600 1.415 0.890 1.460 ;
        RECT 3.115 1.415 3.405 1.460 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dlxtn_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__dlxtn_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__dlxtn_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 1.475 0.955 1.890 1.325 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.330 1.625 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.470 0.785 7.345 1.015 ;
        RECT 0.005 0.105 7.345 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.996000 ;
    PORT
      LAYER li1 ;
        RECT 5.595 1.495 5.895 2.455 ;
        RECT 5.710 1.325 5.895 1.495 ;
        RECT 6.535 1.325 6.805 2.455 ;
        RECT 5.710 0.995 7.235 1.325 ;
        RECT 5.710 0.745 5.895 0.995 ;
        RECT 5.595 0.415 5.895 0.745 ;
        RECT 6.535 0.385 6.805 0.995 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.360 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.895 2.635 ;
        RECT 0.175 1.795 0.890 1.965 ;
        RECT 0.660 0.805 0.890 1.795 ;
        RECT 0.175 0.635 0.890 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.115 0.345 1.285 2.465 ;
        RECT 1.555 1.665 1.885 2.415 ;
        RECT 2.105 1.835 2.420 2.635 ;
        RECT 3.025 2.255 3.950 2.425 ;
        RECT 1.555 1.495 2.290 1.665 ;
        RECT 2.120 1.095 2.290 1.495 ;
        RECT 2.670 1.355 2.955 2.005 ;
        RECT 3.175 1.415 3.565 1.995 ;
        RECT 2.120 0.785 2.540 1.095 ;
        RECT 3.175 1.035 3.345 1.415 ;
        RECT 1.635 0.765 2.540 0.785 ;
        RECT 1.635 0.615 2.290 0.765 ;
        RECT 2.915 0.705 3.345 1.035 ;
        RECT 3.780 1.325 3.950 2.255 ;
        RECT 4.120 2.135 4.290 2.635 ;
        RECT 4.640 1.865 4.860 2.435 ;
        RECT 4.140 1.535 4.860 1.865 ;
        RECT 4.670 1.325 4.860 1.535 ;
        RECT 5.090 1.495 5.375 2.635 ;
        RECT 6.065 1.495 6.315 2.635 ;
        RECT 7.005 1.495 7.175 2.635 ;
        RECT 3.780 0.995 4.500 1.325 ;
        RECT 4.670 0.995 5.490 1.325 ;
        RECT 1.635 0.345 1.805 0.615 ;
        RECT 3.780 0.535 3.950 0.995 ;
        RECT 1.975 0.085 2.355 0.445 ;
        RECT 3.090 0.365 3.950 0.535 ;
        RECT 4.120 0.085 4.290 0.610 ;
        RECT 4.670 0.415 4.860 0.995 ;
        RECT 5.090 0.085 5.375 0.715 ;
        RECT 6.065 0.085 6.315 0.825 ;
        RECT 7.005 0.085 7.175 0.715 ;
        RECT 0.000 -0.085 7.360 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 0.660 1.400 0.830 1.570 ;
        RECT 1.115 1.770 1.285 1.940 ;
        RECT 2.670 1.770 2.840 1.940 ;
        RECT 3.175 1.400 3.345 1.570 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
      LAYER met1 ;
        RECT 1.055 1.940 1.345 1.970 ;
        RECT 2.610 1.940 2.900 1.970 ;
        RECT 1.055 1.800 2.900 1.940 ;
        RECT 1.055 1.740 1.345 1.800 ;
        RECT 2.610 1.740 2.900 1.800 ;
        RECT 0.600 1.460 3.410 1.600 ;
        RECT 0.600 1.370 0.890 1.460 ;
        RECT 3.115 1.370 3.410 1.460 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dlxtn_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__dlygate4sd1_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__dlygate4sd1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.055 0.605 1.615 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.465 0.785 3.200 1.015 ;
        RECT 0.005 0.105 3.200 0.785 ;
        RECT 0.140 -0.085 0.310 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.449000 ;
    PORT
      LAYER li1 ;
        RECT 2.860 1.495 3.120 2.465 ;
        RECT 2.950 0.825 3.120 1.495 ;
        RECT 2.830 0.255 3.120 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.085 2.005 0.380 2.465 ;
        RECT 0.600 2.175 0.815 2.635 ;
        RECT 0.985 2.175 1.420 2.465 ;
        RECT 0.085 1.785 0.945 2.005 ;
        RECT 0.775 1.325 0.945 1.785 ;
        RECT 0.775 0.995 1.080 1.325 ;
        RECT 1.250 1.275 1.420 2.175 ;
        RECT 1.615 1.745 1.840 2.430 ;
        RECT 2.145 1.915 2.515 2.635 ;
        RECT 1.615 1.575 2.610 1.745 ;
        RECT 2.400 1.325 2.610 1.575 ;
        RECT 1.250 1.075 2.000 1.275 ;
        RECT 0.775 0.885 0.945 0.995 ;
        RECT 0.095 0.715 0.945 0.885 ;
        RECT 0.095 0.255 0.380 0.715 ;
        RECT 1.250 0.545 1.420 1.075 ;
        RECT 2.400 0.995 2.730 1.325 ;
        RECT 2.400 0.905 2.610 0.995 ;
        RECT 0.600 0.085 0.815 0.545 ;
        RECT 0.985 0.255 1.420 0.545 ;
        RECT 1.615 0.735 2.610 0.905 ;
        RECT 1.615 0.255 1.840 0.735 ;
        RECT 2.145 0.085 2.555 0.565 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dlygate4sd1_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__dlygate4sd2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__dlygate4sd2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.055 0.605 1.615 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.465 0.785 3.200 1.015 ;
        RECT 0.005 0.105 3.200 0.785 ;
        RECT 0.140 -0.085 0.310 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.464000 ;
    PORT
      LAYER li1 ;
        RECT 2.780 1.495 3.110 2.465 ;
        RECT 2.860 0.825 3.110 1.495 ;
        RECT 2.780 0.255 3.110 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.085 2.005 0.380 2.465 ;
        RECT 0.600 2.175 0.815 2.635 ;
        RECT 0.985 2.175 1.420 2.465 ;
        RECT 0.085 1.785 0.945 2.005 ;
        RECT 0.775 1.325 0.945 1.785 ;
        RECT 0.775 0.995 1.080 1.325 ;
        RECT 1.250 1.275 1.420 2.175 ;
        RECT 1.615 1.745 1.840 2.080 ;
        RECT 2.145 1.915 2.515 2.635 ;
        RECT 1.615 1.575 2.610 1.745 ;
        RECT 2.400 1.325 2.610 1.575 ;
        RECT 1.250 1.075 2.095 1.275 ;
        RECT 0.775 0.885 0.945 0.995 ;
        RECT 0.095 0.715 0.945 0.885 ;
        RECT 0.095 0.255 0.380 0.715 ;
        RECT 1.250 0.545 1.420 1.075 ;
        RECT 2.400 0.995 2.690 1.325 ;
        RECT 2.400 0.905 2.610 0.995 ;
        RECT 0.600 0.085 0.815 0.545 ;
        RECT 0.985 0.255 1.420 0.545 ;
        RECT 1.615 0.735 2.610 0.905 ;
        RECT 1.615 0.510 1.840 0.735 ;
        RECT 2.145 0.085 2.555 0.565 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dlygate4sd2_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__dlygate4sd3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__dlygate4sd3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.055 0.605 1.615 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.765 0.785 3.610 1.015 ;
        RECT 0.005 0.335 3.610 0.785 ;
        RECT 0.005 0.105 1.755 0.335 ;
        RECT 2.600 0.105 3.610 0.335 ;
        RECT 0.140 -0.085 0.310 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 3.190 1.495 3.595 2.465 ;
        RECT 3.325 0.825 3.595 1.495 ;
        RECT 3.190 0.255 3.595 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.085 2.005 0.380 2.465 ;
        RECT 0.605 2.175 0.855 2.635 ;
        RECT 1.305 2.175 1.740 2.465 ;
        RECT 0.085 1.785 0.945 2.005 ;
        RECT 0.775 1.325 0.945 1.785 ;
        RECT 0.775 0.995 1.400 1.325 ;
        RECT 1.570 1.275 1.740 2.175 ;
        RECT 1.910 1.745 2.130 2.080 ;
        RECT 2.690 1.915 3.020 2.635 ;
        RECT 1.910 1.575 3.020 1.745 ;
        RECT 2.810 1.325 3.020 1.575 ;
        RECT 1.570 1.075 2.475 1.275 ;
        RECT 0.775 0.885 0.945 0.995 ;
        RECT 0.095 0.715 0.945 0.885 ;
        RECT 0.095 0.255 0.380 0.715 ;
        RECT 1.570 0.545 1.740 1.075 ;
        RECT 2.810 0.995 3.155 1.325 ;
        RECT 2.810 0.905 3.020 0.995 ;
        RECT 0.600 0.085 0.815 0.545 ;
        RECT 1.305 0.255 1.740 0.545 ;
        RECT 1.910 0.735 3.020 0.905 ;
        RECT 1.910 0.510 2.140 0.735 ;
        RECT 2.690 0.085 3.020 0.565 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dlygate4sd3_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__ebufn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__ebufn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.355 1.615 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.358200 ;
    PORT
      LAYER li1 ;
        RECT 0.960 1.075 1.290 1.630 ;
    END
  END TE_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.540 0.785 3.675 1.015 ;
        RECT 0.005 0.335 3.675 0.785 ;
        RECT 0.005 0.105 1.005 0.335 ;
        RECT 2.175 0.105 3.675 0.335 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.700500 ;
    PORT
      LAYER li1 ;
        RECT 2.125 1.495 3.585 2.465 ;
        RECT 3.315 0.825 3.585 1.495 ;
        RECT 3.255 0.255 3.585 0.825 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT -0.005 2.635 3.680 2.805 ;
        RECT 0.085 2.005 0.345 2.465 ;
        RECT 0.515 2.175 0.890 2.635 ;
        RECT 1.115 2.005 1.370 2.460 ;
        RECT 1.540 2.175 1.900 2.635 ;
        RECT 0.085 1.785 0.790 2.005 ;
        RECT 1.115 1.800 1.905 2.005 ;
        RECT 0.525 0.825 0.790 1.785 ;
        RECT 1.460 1.325 1.905 1.800 ;
        RECT 1.460 1.075 2.745 1.325 ;
        RECT 0.085 0.615 1.235 0.825 ;
        RECT 1.460 0.635 1.790 1.075 ;
        RECT 2.915 0.995 3.145 1.325 ;
        RECT 2.915 0.905 3.085 0.995 ;
        RECT 1.960 0.735 3.085 0.905 ;
        RECT 0.085 0.280 0.345 0.615 ;
        RECT 1.065 0.465 1.235 0.615 ;
        RECT 1.960 0.465 2.175 0.735 ;
        RECT 0.515 0.085 0.895 0.445 ;
        RECT 1.065 0.255 2.175 0.465 ;
        RECT 2.345 0.085 3.085 0.565 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__ebufn_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__ebufn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__ebufn_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.765 0.775 1.675 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.516600 ;
    PORT
      LAYER li1 ;
        RECT 0.945 0.765 1.300 1.275 ;
    END
  END TE_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.930 0.785 4.485 1.015 ;
        RECT 0.005 0.105 4.485 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.530500 ;
    PORT
      LAYER li1 ;
        RECT 3.595 1.765 3.995 2.125 ;
        RECT 1.985 1.625 3.995 1.765 ;
        RECT 1.985 1.445 4.460 1.625 ;
        RECT 4.230 0.855 4.460 1.445 ;
        RECT 3.545 0.635 4.460 0.855 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.085 0.280 0.345 2.465 ;
        RECT 0.515 1.845 1.000 2.635 ;
        RECT 1.220 1.765 1.510 2.465 ;
        RECT 1.700 2.105 1.910 2.465 ;
        RECT 2.080 2.275 2.460 2.635 ;
        RECT 2.680 2.295 4.425 2.465 ;
        RECT 2.680 2.105 3.375 2.295 ;
        RECT 1.700 1.935 3.375 2.105 ;
        RECT 4.165 1.795 4.425 2.295 ;
        RECT 1.220 1.445 1.815 1.765 ;
        RECT 1.550 1.275 1.815 1.445 ;
        RECT 1.550 1.025 3.215 1.275 ;
        RECT 3.495 1.025 3.955 1.275 ;
        RECT 1.550 0.595 1.830 1.025 ;
        RECT 0.515 0.085 0.900 0.595 ;
        RECT 1.070 0.255 1.830 0.595 ;
        RECT 2.000 0.655 3.375 0.855 ;
        RECT 2.000 0.255 2.320 0.655 ;
        RECT 2.490 0.085 2.870 0.485 ;
        RECT 3.090 0.465 3.375 0.655 ;
        RECT 3.090 0.275 4.400 0.465 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.150 1.060 0.320 1.230 ;
        RECT 3.680 1.060 3.850 1.230 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
      LAYER met1 ;
        RECT 0.085 1.120 3.910 1.260 ;
        RECT 0.085 1.030 0.380 1.120 ;
        RECT 3.570 1.030 3.910 1.120 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__ebufn_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__ebufn_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__ebufn_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.490 0.765 0.830 1.675 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.954300 ;
    PORT
      LAYER li1 ;
        RECT 1.000 0.765 1.380 1.425 ;
    END
  END TE_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 6.395 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.028500 ;
    PORT
      LAYER li1 ;
        RECT 1.995 1.445 6.335 1.725 ;
        RECT 6.105 0.855 6.335 1.445 ;
        RECT 4.495 0.615 6.335 0.855 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.085 1.765 0.345 2.465 ;
        RECT 0.515 1.845 0.980 2.635 ;
        RECT 1.200 1.765 1.455 2.465 ;
        RECT 1.665 2.105 1.910 2.465 ;
        RECT 2.080 2.275 2.460 2.635 ;
        RECT 2.680 2.105 2.850 2.465 ;
        RECT 3.070 2.275 3.400 2.635 ;
        RECT 3.620 2.105 6.285 2.465 ;
        RECT 1.665 1.935 6.285 2.105 ;
        RECT 1.995 1.895 6.285 1.935 ;
        RECT 0.085 0.665 0.320 1.765 ;
        RECT 1.200 1.595 1.825 1.765 ;
        RECT 1.550 1.275 1.825 1.595 ;
        RECT 1.550 1.025 4.160 1.275 ;
        RECT 4.330 1.025 5.935 1.275 ;
        RECT 0.085 0.280 0.345 0.665 ;
        RECT 1.550 0.595 1.825 1.025 ;
        RECT 0.515 0.085 0.980 0.595 ;
        RECT 1.200 0.255 1.825 0.595 ;
        RECT 1.995 0.655 4.325 0.855 ;
        RECT 1.995 0.255 2.325 0.655 ;
        RECT 2.495 0.085 2.875 0.485 ;
        RECT 3.095 0.275 3.265 0.655 ;
        RECT 3.435 0.085 3.815 0.485 ;
        RECT 4.035 0.445 4.325 0.655 ;
        RECT 4.035 0.255 6.285 0.445 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.150 1.105 0.320 1.275 ;
        RECT 4.710 1.105 4.880 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
      LAYER met1 ;
        RECT 0.085 1.165 4.940 1.305 ;
        RECT 0.085 1.075 0.380 1.165 ;
        RECT 4.650 1.075 4.940 1.165 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__ebufn_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__ebufn_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__ebufn_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.040 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.430 1.615 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.631100 ;
    PORT
      LAYER li1 ;
        RECT 1.020 1.325 1.405 1.695 ;
        RECT 1.020 0.995 1.530 1.325 ;
        RECT 1.020 0.620 1.405 0.995 ;
    END
  END TE_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.040 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 11.005 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 11.230 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.040 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.024500 ;
    PORT
      LAYER li1 ;
        RECT 2.145 1.445 10.925 1.725 ;
        RECT 10.675 0.855 10.925 1.445 ;
        RECT 7.225 0.615 10.925 0.855 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 11.040 2.805 ;
        RECT 0.085 1.785 0.445 2.635 ;
        RECT 0.665 1.615 0.850 2.465 ;
        RECT 1.020 1.865 1.405 2.635 ;
        RECT 0.085 0.085 0.445 0.825 ;
        RECT 0.650 0.280 0.850 1.615 ;
        RECT 1.575 1.495 1.975 2.465 ;
        RECT 2.145 2.065 2.395 2.465 ;
        RECT 2.565 2.235 2.995 2.635 ;
        RECT 3.215 2.065 3.385 2.465 ;
        RECT 3.605 2.235 4.035 2.635 ;
        RECT 4.255 2.065 4.425 2.465 ;
        RECT 4.645 2.235 5.075 2.635 ;
        RECT 5.295 2.065 5.465 2.465 ;
        RECT 5.685 2.235 6.115 2.635 ;
        RECT 6.335 2.065 10.925 2.465 ;
        RECT 2.145 1.895 10.925 2.065 ;
        RECT 1.750 1.275 1.975 1.495 ;
        RECT 1.750 1.025 6.875 1.275 ;
        RECT 7.125 1.025 10.455 1.275 ;
        RECT 1.750 0.825 2.135 1.025 ;
        RECT 1.020 0.085 1.405 0.445 ;
        RECT 1.575 0.255 2.135 0.825 ;
        RECT 2.305 0.655 7.055 0.855 ;
        RECT 2.305 0.255 2.685 0.655 ;
        RECT 2.855 0.085 3.285 0.485 ;
        RECT 3.505 0.275 3.725 0.655 ;
        RECT 3.895 0.085 4.325 0.485 ;
        RECT 4.545 0.255 4.765 0.655 ;
        RECT 4.935 0.085 5.365 0.485 ;
        RECT 5.585 0.275 5.805 0.655 ;
        RECT 5.975 0.085 6.405 0.485 ;
        RECT 6.625 0.445 7.055 0.655 ;
        RECT 6.625 0.255 10.925 0.445 ;
        RECT 0.000 -0.085 11.040 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 0.655 1.060 0.825 1.230 ;
        RECT 7.630 1.060 7.800 1.230 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
      LAYER met1 ;
        RECT 0.545 1.120 7.860 1.260 ;
        RECT 0.545 1.030 0.885 1.120 ;
        RECT 7.520 1.030 7.860 1.120 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__ebufn_8

#--------EOF---------

MACRO sky130_fd_sc_hdll__einvn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__einvn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.430 0.765 2.675 1.615 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.358200 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.955 0.510 1.725 ;
    END
  END TE_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.540 0.785 2.755 1.015 ;
        RECT 0.005 0.105 2.755 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.471500 ;
    PORT
      LAYER li1 ;
        RECT 1.400 1.785 2.675 2.465 ;
        RECT 1.970 0.595 2.210 1.785 ;
        RECT 1.970 0.255 2.675 0.595 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.085 2.065 0.370 2.465 ;
        RECT 0.540 2.235 0.920 2.635 ;
        RECT 0.085 1.895 0.920 2.065 ;
        RECT 0.735 1.615 0.920 1.895 ;
        RECT 0.735 1.440 1.600 1.615 ;
        RECT 1.120 0.805 1.600 1.440 ;
        RECT 0.735 0.785 1.600 0.805 ;
        RECT 0.085 0.615 1.600 0.785 ;
        RECT 0.085 0.255 0.370 0.615 ;
        RECT 0.540 0.085 1.590 0.445 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__einvn_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__einvn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__einvn_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.985 1.075 3.535 1.275 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.516600 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.325 1.385 ;
    END
  END TE_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.040 0.785 3.505 1.015 ;
        RECT 0.005 0.105 3.505 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.768000 ;
    PORT
      LAYER li1 ;
        RECT 3.035 1.695 3.535 2.465 ;
        RECT 2.145 1.445 3.535 1.695 ;
        RECT 2.445 0.595 2.815 1.445 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.085 1.725 0.345 2.465 ;
        RECT 0.515 1.895 0.945 2.635 ;
        RECT 1.170 2.085 1.340 2.465 ;
        RECT 1.510 2.255 2.475 2.635 ;
        RECT 2.695 2.085 2.865 2.465 ;
        RECT 1.170 1.865 2.865 2.085 ;
        RECT 0.085 1.555 0.945 1.725 ;
        RECT 0.495 1.275 0.945 1.555 ;
        RECT 1.170 1.445 1.925 1.865 ;
        RECT 0.495 0.995 2.180 1.275 ;
        RECT 0.495 0.825 0.890 0.995 ;
        RECT 0.085 0.655 0.890 0.825 ;
        RECT 1.065 0.655 2.270 0.825 ;
        RECT 0.085 0.255 0.345 0.655 ;
        RECT 0.515 0.085 0.895 0.485 ;
        RECT 1.065 0.255 1.380 0.655 ;
        RECT 1.600 0.085 1.930 0.485 ;
        RECT 2.100 0.425 2.270 0.655 ;
        RECT 3.165 0.425 3.435 0.775 ;
        RECT 2.100 0.255 3.435 0.425 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__einvn_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__einvn_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__einvn_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 4.980 0.620 5.415 1.325 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.954300 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.345 1.325 ;
    END
  END TE_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.390 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.996000 ;
    PORT
      LAYER li1 ;
        RECT 3.490 1.480 3.870 2.075 ;
        RECT 4.430 1.480 4.810 2.075 ;
        RECT 3.490 0.620 4.810 1.480 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.085 1.665 0.345 2.465 ;
        RECT 0.515 1.835 0.895 2.635 ;
        RECT 1.065 1.665 1.340 2.465 ;
        RECT 1.510 1.835 1.890 2.635 ;
        RECT 2.110 1.665 2.280 2.465 ;
        RECT 2.450 1.835 2.890 2.635 ;
        RECT 3.110 2.295 5.200 2.465 ;
        RECT 3.110 1.665 3.320 2.295 ;
        RECT 0.085 1.495 0.895 1.665 ;
        RECT 1.065 1.495 3.320 1.665 ;
        RECT 4.090 1.650 4.260 2.295 ;
        RECT 5.030 1.650 5.200 2.295 ;
        RECT 0.515 1.325 0.895 1.495 ;
        RECT 0.515 0.995 3.320 1.325 ;
        RECT 0.515 0.825 0.895 0.995 ;
        RECT 0.085 0.655 0.895 0.825 ;
        RECT 1.065 0.655 3.295 0.825 ;
        RECT 0.085 0.255 0.345 0.655 ;
        RECT 0.515 0.085 0.895 0.485 ;
        RECT 1.065 0.255 1.385 0.655 ;
        RECT 1.605 0.085 1.935 0.485 ;
        RECT 2.155 0.255 2.325 0.655 ;
        RECT 2.545 0.085 2.875 0.485 ;
        RECT 3.125 0.450 3.295 0.655 ;
        RECT 3.125 0.255 5.435 0.450 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__einvn_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__einvn_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__einvn_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.200 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.220000 ;
    PORT
      LAYER li1 ;
        RECT 5.145 0.995 8.650 1.285 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.631100 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.995 0.345 1.325 ;
    END
  END TE_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.200 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 9.150 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.390 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.200 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.024500 ;
    PORT
      LAYER li1 ;
        RECT 5.370 1.625 5.750 2.125 ;
        RECT 6.310 1.625 6.690 2.125 ;
        RECT 7.250 1.625 7.630 2.125 ;
        RECT 8.190 1.625 8.570 2.125 ;
        RECT 5.370 1.455 9.095 1.625 ;
        RECT 8.870 0.825 9.095 1.455 ;
        RECT 5.370 0.620 9.095 0.825 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.200 2.805 ;
        RECT 0.090 1.665 0.345 2.465 ;
        RECT 0.515 1.835 0.895 2.635 ;
        RECT 1.065 1.665 1.340 2.465 ;
        RECT 1.510 1.835 1.890 2.635 ;
        RECT 2.110 1.665 2.280 2.465 ;
        RECT 2.450 1.835 2.830 2.635 ;
        RECT 3.050 1.665 3.220 2.465 ;
        RECT 3.390 1.835 3.770 2.635 ;
        RECT 3.990 1.665 4.160 2.465 ;
        RECT 4.330 1.835 4.730 2.635 ;
        RECT 4.950 2.295 9.095 2.465 ;
        RECT 4.950 1.665 5.200 2.295 ;
        RECT 5.970 1.795 6.140 2.295 ;
        RECT 6.910 1.795 7.080 2.295 ;
        RECT 7.850 1.795 8.020 2.295 ;
        RECT 8.790 1.795 9.095 2.295 ;
        RECT 0.090 1.495 0.895 1.665 ;
        RECT 1.065 1.495 5.200 1.665 ;
        RECT 0.515 1.325 0.895 1.495 ;
        RECT 0.515 0.995 4.975 1.325 ;
        RECT 0.515 0.825 0.895 0.995 ;
        RECT 0.090 0.655 0.895 0.825 ;
        RECT 1.065 0.655 5.200 0.825 ;
        RECT 0.090 0.255 0.345 0.655 ;
        RECT 0.515 0.085 0.895 0.485 ;
        RECT 1.065 0.255 1.385 0.655 ;
        RECT 1.605 0.085 1.935 0.485 ;
        RECT 2.155 0.255 2.325 0.655 ;
        RECT 2.545 0.085 2.875 0.485 ;
        RECT 3.095 0.255 3.265 0.655 ;
        RECT 3.485 0.085 3.815 0.485 ;
        RECT 4.035 0.255 4.205 0.655 ;
        RECT 4.425 0.085 4.765 0.485 ;
        RECT 4.985 0.450 5.200 0.655 ;
        RECT 4.985 0.255 9.095 0.450 ;
        RECT 0.000 -0.085 9.200 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__einvn_8

#--------EOF---------

MACRO sky130_fd_sc_hdll__einvp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__einvp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.385 0.975 2.625 1.955 ;
    END
  END A
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.236100 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.595 1.725 ;
    END
  END TE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.490 0.785 2.705 1.015 ;
        RECT 0.005 0.105 2.705 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.488000 ;
    PORT
      LAYER li1 ;
        RECT 1.980 2.125 2.625 2.465 ;
        RECT 1.980 0.805 2.155 2.125 ;
        RECT 1.980 0.255 2.625 0.805 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.085 2.065 0.345 2.465 ;
        RECT 0.515 2.235 1.740 2.635 ;
        RECT 0.085 1.895 1.690 2.065 ;
        RECT 0.765 0.825 1.690 1.895 ;
        RECT 0.085 0.655 1.690 0.825 ;
        RECT 0.085 0.255 0.345 0.655 ;
        RECT 0.515 0.085 1.500 0.485 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__einvp_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__einvp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__einvp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 3.245 0.765 3.535 1.615 ;
    END
  END A
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373200 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.330 1.615 ;
    END
  END TE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.540 0.785 3.585 1.015 ;
        RECT 0.005 0.105 3.585 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.530500 ;
    PORT
      LAYER li1 ;
        RECT 2.645 0.595 3.075 2.125 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.085 1.955 0.345 2.465 ;
        RECT 0.515 2.125 0.925 2.635 ;
        RECT 0.085 1.785 0.925 1.955 ;
        RECT 0.500 1.325 0.925 1.785 ;
        RECT 1.145 1.725 1.385 2.465 ;
        RECT 1.605 1.895 1.935 2.635 ;
        RECT 2.185 2.295 3.530 2.465 ;
        RECT 2.185 1.725 2.355 2.295 ;
        RECT 3.245 1.785 3.530 2.295 ;
        RECT 1.145 1.555 2.355 1.725 ;
        RECT 0.500 0.995 2.105 1.325 ;
        RECT 0.500 0.825 0.925 0.995 ;
        RECT 0.085 0.655 0.925 0.825 ;
        RECT 1.145 0.655 2.475 0.825 ;
        RECT 0.085 0.255 0.345 0.655 ;
        RECT 0.515 0.085 0.925 0.485 ;
        RECT 1.145 0.255 1.340 0.655 ;
        RECT 1.510 0.085 1.880 0.485 ;
        RECT 2.140 0.425 2.475 0.655 ;
        RECT 3.245 0.425 3.530 0.595 ;
        RECT 2.140 0.255 3.530 0.425 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__einvp_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__einvp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__einvp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 4.210 1.020 5.410 1.275 ;
    END
  END A
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.667500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.330 1.615 ;
    END
  END TE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.390 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.996000 ;
    PORT
      LAYER li1 ;
        RECT 3.490 1.615 3.870 2.125 ;
        RECT 4.430 1.615 4.810 2.125 ;
        RECT 3.490 1.445 4.810 1.615 ;
        RECT 3.490 0.850 4.030 1.445 ;
        RECT 3.490 0.635 5.410 0.850 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.085 1.955 0.345 2.465 ;
        RECT 0.515 2.125 0.925 2.635 ;
        RECT 0.085 1.785 0.925 1.955 ;
        RECT 0.500 1.325 0.925 1.785 ;
        RECT 1.175 1.725 1.385 2.465 ;
        RECT 1.605 1.895 1.935 2.635 ;
        RECT 2.155 1.725 2.325 2.465 ;
        RECT 2.545 1.895 2.905 2.635 ;
        RECT 3.125 2.295 5.410 2.465 ;
        RECT 3.125 1.725 3.295 2.295 ;
        RECT 4.090 1.785 4.260 2.295 ;
        RECT 1.175 1.555 3.295 1.725 ;
        RECT 5.030 1.445 5.410 2.295 ;
        RECT 0.500 0.995 3.320 1.325 ;
        RECT 0.500 0.825 0.745 0.995 ;
        RECT 0.085 0.655 0.745 0.825 ;
        RECT 1.135 0.655 3.320 0.825 ;
        RECT 0.085 0.255 0.345 0.655 ;
        RECT 0.515 0.085 0.895 0.485 ;
        RECT 1.135 0.255 1.305 0.655 ;
        RECT 1.475 0.085 1.855 0.485 ;
        RECT 2.075 0.255 2.245 0.655 ;
        RECT 2.415 0.085 2.805 0.485 ;
        RECT 2.985 0.465 3.320 0.655 ;
        RECT 2.985 0.255 5.410 0.465 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__einvp_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__einvp_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__einvp_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.200 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.220000 ;
    PORT
      LAYER li1 ;
        RECT 6.020 1.020 9.050 1.275 ;
    END
  END A
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.330 1.615 ;
    END
  END TE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.200 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 9.150 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.390 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.200 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.992000 ;
    PORT
      LAYER li1 ;
        RECT 5.370 1.615 5.750 2.125 ;
        RECT 6.310 1.615 6.690 2.125 ;
        RECT 7.250 1.615 7.630 2.125 ;
        RECT 8.190 1.615 8.570 2.125 ;
        RECT 5.370 1.445 8.570 1.615 ;
        RECT 5.370 0.850 5.800 1.445 ;
        RECT 5.370 0.635 9.095 0.850 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.200 2.805 ;
        RECT 0.085 1.955 0.345 2.465 ;
        RECT 0.515 2.125 0.925 2.635 ;
        RECT 0.085 1.785 0.925 1.955 ;
        RECT 0.500 1.325 0.925 1.785 ;
        RECT 1.175 1.725 1.385 2.465 ;
        RECT 1.605 1.895 1.935 2.635 ;
        RECT 2.155 1.725 2.325 2.465 ;
        RECT 2.545 1.895 2.875 2.635 ;
        RECT 3.095 1.725 3.265 2.465 ;
        RECT 3.485 1.895 3.815 2.635 ;
        RECT 4.035 1.725 4.205 2.465 ;
        RECT 4.425 1.895 4.755 2.635 ;
        RECT 4.975 2.295 9.095 2.465 ;
        RECT 4.975 1.725 5.200 2.295 ;
        RECT 5.970 1.785 6.140 2.295 ;
        RECT 6.910 1.785 7.080 2.295 ;
        RECT 7.850 1.785 8.020 2.295 ;
        RECT 1.175 1.555 5.200 1.725 ;
        RECT 8.790 1.445 9.095 2.295 ;
        RECT 0.500 0.995 5.200 1.325 ;
        RECT 0.500 0.825 0.745 0.995 ;
        RECT 0.085 0.655 0.745 0.825 ;
        RECT 1.135 0.655 5.200 0.825 ;
        RECT 0.085 0.255 0.345 0.655 ;
        RECT 0.515 0.085 0.895 0.485 ;
        RECT 1.135 0.255 1.305 0.655 ;
        RECT 1.475 0.085 1.855 0.485 ;
        RECT 2.075 0.255 2.245 0.655 ;
        RECT 2.415 0.085 2.795 0.485 ;
        RECT 3.015 0.255 3.185 0.655 ;
        RECT 3.355 0.085 3.735 0.485 ;
        RECT 3.955 0.255 4.125 0.655 ;
        RECT 4.295 0.085 4.685 0.485 ;
        RECT 4.855 0.465 5.200 0.655 ;
        RECT 4.855 0.255 9.095 0.465 ;
        RECT 0.000 -0.085 9.200 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__einvp_8

#--------EOF---------

MACRO sky130_fd_sc_hdll__fill_1
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hdll__fill_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.460 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 0.460 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.140 -0.055 0.260 0.055 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 0.650 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 0.460 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 0.460 2.805 ;
        RECT 0.000 -0.085 0.460 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__fill_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__fill_2
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hdll__fill_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.920 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 0.920 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.155 -0.050 0.315 0.060 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 1.110 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 0.920 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 0.920 2.805 ;
        RECT 0.000 -0.085 0.920 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__fill_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__fill_4
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hdll__fill_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.175 -0.060 0.285 0.060 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.840 2.805 ;
        RECT 0.000 -0.085 1.840 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__fill_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__fill_8
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hdll__fill_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.130 -0.120 0.350 0.050 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__fill_8

#--------EOF---------

MACRO sky130_fd_sc_hdll__inputiso0n_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__inputiso0n_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.100 1.325 0.365 1.685 ;
        RECT 0.100 1.075 0.590 1.325 ;
    END
  END A
  PIN SLEEP_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.855 1.075 1.275 1.325 ;
    END
  END SLEEP_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.085 0.925 2.015 1.015 ;
        RECT 0.005 0.245 2.015 0.925 ;
        RECT 0.145 0.105 2.015 0.245 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.539000 ;
    PORT
      LAYER li1 ;
        RECT 1.745 1.915 2.205 2.465 ;
        RECT 1.955 0.545 2.205 1.915 ;
        RECT 1.595 0.255 2.205 0.545 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.125 1.965 0.405 2.635 ;
        RECT 0.625 1.745 0.925 2.295 ;
        RECT 1.175 1.915 1.505 2.635 ;
        RECT 0.625 1.575 1.695 1.745 ;
        RECT 1.525 0.905 1.695 1.575 ;
        RECT 0.125 0.715 1.695 0.905 ;
        RECT 0.125 0.355 0.455 0.715 ;
        RECT 1.175 0.085 1.425 0.545 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__inputiso0n_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__inputiso0p_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__inputiso0p_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.645 1.835 1.955 ;
    END
  END A
  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.765 0.445 1.615 ;
    END
  END SLEEP
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.990 0.785 2.960 1.015 ;
        RECT 0.005 0.105 2.960 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 2.505 1.580 3.080 2.365 ;
        RECT 2.905 0.775 3.080 1.580 ;
        RECT 2.620 0.255 3.080 0.775 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.175 2.015 0.345 2.445 ;
        RECT 0.515 2.185 0.895 2.635 ;
        RECT 0.175 1.785 0.895 2.015 ;
        RECT 0.645 1.135 0.895 1.785 ;
        RECT 1.065 1.475 1.335 2.420 ;
        RECT 1.565 2.165 2.325 2.635 ;
        RECT 1.065 1.325 1.885 1.475 ;
        RECT 1.065 1.305 2.475 1.325 ;
        RECT 0.645 0.805 1.180 1.135 ;
        RECT 1.350 0.945 2.475 1.305 ;
        RECT 0.090 0.085 0.425 0.590 ;
        RECT 0.645 0.280 0.885 0.805 ;
        RECT 1.350 0.610 1.590 0.945 ;
        RECT 1.165 0.415 1.590 0.610 ;
        RECT 1.165 0.270 1.335 0.415 ;
        RECT 2.070 0.085 2.400 0.580 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__inputiso0p_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__inputiso1n_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__inputiso1n_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.540 2.085 1.895 2.415 ;
    END
  END A
  PIN SLEEP_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 0.425 1.325 ;
    END
  END SLEEP_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.020 0.815 3.025 1.015 ;
        RECT 0.005 0.135 3.025 0.815 ;
        RECT 0.150 -0.085 0.320 0.135 ;
        RECT 2.020 0.105 3.025 0.135 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.472000 ;
    PORT
      LAYER li1 ;
        RECT 2.675 1.495 3.080 2.465 ;
        RECT 2.910 0.760 3.080 1.495 ;
        RECT 2.675 0.415 3.080 0.760 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.090 1.495 0.345 2.635 ;
        RECT 0.645 1.325 0.815 1.885 ;
        RECT 1.040 1.665 1.460 1.915 ;
        RECT 2.125 1.835 2.405 2.635 ;
        RECT 1.040 1.495 2.505 1.665 ;
        RECT 0.645 0.995 1.385 1.325 ;
        RECT 0.645 0.905 0.895 0.995 ;
        RECT 0.110 0.735 0.895 0.905 ;
        RECT 2.335 0.825 2.505 1.495 ;
        RECT 0.110 0.265 0.420 0.735 ;
        RECT 1.655 0.655 2.505 0.825 ;
        RECT 0.640 0.085 1.375 0.565 ;
        RECT 1.655 0.305 1.825 0.655 ;
        RECT 1.995 0.085 2.425 0.485 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__inputiso1n_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__inputiso1p_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__inputiso1p_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.440 1.325 ;
    END
  END A
  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.000 0.765 1.315 1.325 ;
    END
  END SLEEP
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.095 0.785 2.135 1.015 ;
        RECT 0.090 0.105 2.135 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.650500 ;
    PORT
      LAYER li1 ;
        RECT 1.795 1.845 2.215 2.465 ;
        RECT 1.900 0.825 2.215 1.845 ;
        RECT 1.665 0.255 2.215 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.150 1.665 0.540 1.840 ;
        RECT 1.185 1.835 1.515 2.635 ;
        RECT 0.150 1.495 1.705 1.665 ;
        RECT 0.610 0.595 0.830 1.495 ;
        RECT 1.535 0.995 1.705 1.495 ;
        RECT 0.190 0.085 0.430 0.595 ;
        RECT 0.610 0.265 0.940 0.595 ;
        RECT 1.220 0.085 1.435 0.595 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__inputiso1p_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__inv_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__inv_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.075 0.650 1.315 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.210 0.105 1.190 1.015 ;
        RECT 0.210 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 1.570 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 0.770 1.485 1.285 2.465 ;
        RECT 0.995 0.885 1.285 1.485 ;
        RECT 0.770 0.255 1.285 0.885 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.380 2.805 ;
        RECT 0.340 1.495 0.550 2.635 ;
        RECT 0.320 0.085 0.550 0.905 ;
        RECT 0.000 -0.085 1.380 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__inv_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__inv_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__inv_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 0.435 1.325 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.015 0.105 1.465 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.498000 ;
    PORT
      LAYER li1 ;
        RECT 0.525 1.485 0.905 2.465 ;
        RECT 0.605 0.885 0.905 1.485 ;
        RECT 0.525 0.255 0.905 0.885 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.840 2.805 ;
        RECT 0.125 1.495 0.355 2.635 ;
        RECT 1.125 1.495 1.335 2.635 ;
        RECT 0.125 0.085 0.355 0.905 ;
        RECT 1.125 0.085 1.335 0.905 ;
        RECT 0.000 -0.085 1.840 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__inv_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__inv_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__inv_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 1.885 1.325 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.055 0.105 2.690 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.996000 ;
    PORT
      LAYER li1 ;
        RECT 0.565 1.665 0.945 2.465 ;
        RECT 1.505 1.685 1.885 2.465 ;
        RECT 1.505 1.665 2.665 1.685 ;
        RECT 0.565 1.495 2.665 1.665 ;
        RECT 2.395 0.905 2.665 1.495 ;
        RECT 0.565 0.725 2.665 0.905 ;
        RECT 0.565 0.255 0.945 0.725 ;
        RECT 1.505 0.255 1.885 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.130 1.495 0.395 2.635 ;
        RECT 1.165 1.835 1.335 2.635 ;
        RECT 2.105 2.175 2.315 2.635 ;
        RECT 0.130 0.085 0.395 0.545 ;
        RECT 1.165 0.085 1.335 0.545 ;
        RECT 2.105 0.085 2.355 0.550 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__inv_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__inv_6
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__inv_6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.665000 ;
    PORT
      LAYER li1 ;
        RECT 0.285 1.075 2.695 1.325 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.055 0.105 3.345 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.494000 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.665 0.895 2.465 ;
        RECT 1.455 1.665 1.835 2.465 ;
        RECT 2.395 1.685 2.775 2.465 ;
        RECT 2.395 1.665 3.265 1.685 ;
        RECT 0.515 1.495 3.265 1.665 ;
        RECT 2.865 0.905 3.265 1.495 ;
        RECT 0.645 0.725 3.265 0.905 ;
        RECT 0.645 0.255 0.815 0.725 ;
        RECT 1.585 0.255 1.755 0.725 ;
        RECT 2.525 0.255 2.695 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.175 1.495 0.345 2.635 ;
        RECT 1.115 1.835 1.285 2.635 ;
        RECT 2.055 1.835 2.225 2.635 ;
        RECT 2.995 2.175 3.165 2.635 ;
        RECT 0.130 0.085 0.395 0.545 ;
        RECT 1.115 0.085 1.285 0.545 ;
        RECT 2.055 0.085 2.225 0.545 ;
        RECT 2.865 0.085 3.165 0.550 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__inv_6

#--------EOF---------

MACRO sky130_fd_sc_hdll__inv_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__inv_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.220000 ;
    PORT
      LAYER li1 ;
        RECT 0.680 1.075 3.885 1.325 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.170 0.105 4.440 1.015 ;
        RECT 0.170 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.024500 ;
    PORT
      LAYER li1 ;
        RECT 0.680 1.665 1.060 2.465 ;
        RECT 1.620 1.665 2.000 2.465 ;
        RECT 2.560 1.665 2.940 2.465 ;
        RECT 3.500 1.665 3.880 2.465 ;
        RECT 0.085 1.495 4.505 1.665 ;
        RECT 0.085 0.905 0.430 1.495 ;
        RECT 4.185 0.905 4.505 1.495 ;
        RECT 0.085 0.715 4.505 0.905 ;
        RECT 0.680 0.255 1.060 0.715 ;
        RECT 1.620 0.255 2.000 0.715 ;
        RECT 2.560 0.255 2.940 0.715 ;
        RECT 3.500 0.255 3.880 0.715 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.255 1.835 0.510 2.635 ;
        RECT 1.280 1.835 1.450 2.635 ;
        RECT 2.220 1.835 2.390 2.635 ;
        RECT 3.160 1.835 3.330 2.635 ;
        RECT 4.100 1.835 4.400 2.635 ;
        RECT 0.255 0.085 0.510 0.545 ;
        RECT 1.280 0.085 1.450 0.545 ;
        RECT 2.220 0.085 2.390 0.545 ;
        RECT 3.160 0.085 3.330 0.545 ;
        RECT 4.100 0.085 4.405 0.545 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__inv_8

#--------EOF---------

MACRO sky130_fd_sc_hdll__inv_12
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__inv_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.330000 ;
    PORT
      LAYER li1 ;
        RECT 0.680 1.075 5.800 1.325 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.170 0.105 6.330 1.015 ;
        RECT 0.170 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.020500 ;
    PORT
      LAYER li1 ;
        RECT 0.680 1.665 1.060 2.465 ;
        RECT 1.620 1.665 2.000 2.465 ;
        RECT 2.560 1.665 2.940 2.465 ;
        RECT 3.500 1.665 3.880 2.465 ;
        RECT 4.440 1.665 4.820 2.465 ;
        RECT 5.380 1.665 5.760 2.465 ;
        RECT 0.085 1.495 6.320 1.665 ;
        RECT 0.085 0.905 0.510 1.495 ;
        RECT 5.970 0.905 6.320 1.495 ;
        RECT 0.085 0.715 6.320 0.905 ;
        RECT 0.680 0.255 1.060 0.715 ;
        RECT 1.620 0.255 2.000 0.715 ;
        RECT 2.560 0.255 2.940 0.715 ;
        RECT 3.500 0.255 3.880 0.715 ;
        RECT 4.440 0.255 4.820 0.715 ;
        RECT 5.380 0.255 5.760 0.715 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.255 1.835 0.510 2.635 ;
        RECT 1.280 1.835 1.450 2.635 ;
        RECT 2.220 1.835 2.390 2.635 ;
        RECT 3.160 1.835 3.330 2.635 ;
        RECT 4.100 1.835 4.270 2.635 ;
        RECT 5.040 1.835 5.210 2.635 ;
        RECT 5.975 1.835 6.230 2.635 ;
        RECT 0.255 0.085 0.510 0.545 ;
        RECT 1.280 0.085 1.450 0.545 ;
        RECT 2.220 0.085 2.390 0.545 ;
        RECT 3.160 0.085 3.330 0.545 ;
        RECT 4.100 0.085 4.270 0.545 ;
        RECT 5.040 0.085 5.210 0.545 ;
        RECT 5.960 0.085 6.230 0.545 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__inv_12

#--------EOF---------

MACRO sky130_fd_sc_hdll__inv_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__inv_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.280 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.440000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 6.125 1.315 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.280 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.070 0.105 8.100 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.470 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.280 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.984000 ;
    PORT
      LAYER li1 ;
        RECT 0.580 1.665 0.960 2.465 ;
        RECT 1.520 1.665 1.900 2.465 ;
        RECT 2.460 1.665 2.840 2.465 ;
        RECT 3.400 1.665 3.780 2.465 ;
        RECT 4.340 1.665 4.720 2.465 ;
        RECT 5.280 1.665 5.660 2.465 ;
        RECT 6.220 1.665 6.600 2.465 ;
        RECT 7.160 1.665 7.540 2.465 ;
        RECT 0.580 1.495 7.540 1.665 ;
        RECT 7.015 0.905 7.540 1.495 ;
        RECT 0.580 0.715 7.540 0.905 ;
        RECT 0.580 0.255 0.960 0.715 ;
        RECT 1.520 0.255 1.900 0.715 ;
        RECT 2.460 0.255 2.840 0.715 ;
        RECT 3.400 0.255 3.780 0.715 ;
        RECT 4.340 0.255 4.720 0.715 ;
        RECT 5.280 0.255 5.660 0.715 ;
        RECT 6.220 0.255 6.600 0.715 ;
        RECT 7.160 0.255 7.540 0.715 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.280 2.805 ;
        RECT 0.200 1.485 0.410 2.635 ;
        RECT 1.180 1.835 1.350 2.635 ;
        RECT 2.120 1.835 2.290 2.635 ;
        RECT 3.060 1.835 3.230 2.635 ;
        RECT 4.000 1.835 4.170 2.635 ;
        RECT 4.940 1.835 5.110 2.635 ;
        RECT 5.880 1.835 6.050 2.635 ;
        RECT 6.820 1.835 6.990 2.635 ;
        RECT 7.760 1.835 7.970 2.635 ;
        RECT 0.180 0.085 0.410 0.885 ;
        RECT 1.180 0.085 1.350 0.545 ;
        RECT 2.120 0.085 2.290 0.545 ;
        RECT 3.060 0.085 3.230 0.545 ;
        RECT 4.000 0.085 4.170 0.545 ;
        RECT 4.940 0.085 5.110 0.545 ;
        RECT 5.880 0.085 6.050 0.545 ;
        RECT 6.820 0.085 6.990 0.545 ;
        RECT 7.760 0.085 7.970 0.885 ;
        RECT 0.000 -0.085 8.280 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__inv_16

#--------EOF---------

MACRO sky130_fd_sc_hdll__isobufsrc_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__isobufsrc_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.100 0.725 0.325 1.325 ;
    END
  END A
  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.010 1.065 1.425 1.325 ;
    END
  END SLEEP
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.775 0.785 2.225 1.015 ;
        RECT 0.240 0.105 2.225 0.785 ;
        RECT 0.240 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.478000 ;
    PORT
      LAYER li1 ;
        RECT 1.755 1.850 2.205 2.465 ;
        RECT 2.025 0.815 2.205 1.850 ;
        RECT 1.285 0.645 2.205 0.815 ;
        RECT 1.285 0.255 1.635 0.645 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.415 1.680 0.675 1.905 ;
        RECT 0.925 1.855 1.255 2.635 ;
        RECT 0.415 1.510 1.855 1.680 ;
        RECT 0.495 0.545 0.675 1.510 ;
        RECT 1.635 0.985 1.855 1.510 ;
        RECT 0.330 0.370 0.675 0.545 ;
        RECT 0.905 0.085 1.115 0.895 ;
        RECT 1.805 0.085 2.135 0.475 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__isobufsrc_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__isobufsrc_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__isobufsrc_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 3.340 1.275 3.555 1.965 ;
        RECT 2.800 1.065 3.555 1.275 ;
    END
  END A
  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.480 1.065 0.970 1.275 ;
    END
  END SLEEP
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.335 3.405 1.015 ;
        RECT 0.010 0.105 2.415 0.335 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.771000 ;
    PORT
      LAYER li1 ;
        RECT 1.525 0.895 1.815 2.125 ;
        RECT 0.535 0.725 1.855 0.895 ;
        RECT 0.535 0.255 0.915 0.725 ;
        RECT 1.475 0.255 1.855 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.085 1.655 0.405 2.465 ;
        RECT 0.625 1.825 0.875 2.635 ;
        RECT 1.095 2.295 2.325 2.465 ;
        RECT 1.095 1.655 1.345 2.295 ;
        RECT 0.085 1.445 1.345 1.655 ;
        RECT 2.035 1.890 2.325 2.295 ;
        RECT 2.035 1.445 2.290 1.890 ;
        RECT 2.595 1.615 2.765 2.460 ;
        RECT 3.025 2.145 3.275 2.635 ;
        RECT 2.460 1.445 2.765 1.615 ;
        RECT 2.460 1.245 2.630 1.445 ;
        RECT 2.075 1.075 2.630 1.245 ;
        RECT 2.415 0.895 2.630 1.075 ;
        RECT 0.085 0.085 0.365 0.895 ;
        RECT 1.135 0.085 1.305 0.555 ;
        RECT 2.075 0.085 2.245 0.895 ;
        RECT 2.415 0.725 2.765 0.895 ;
        RECT 2.595 0.445 2.765 0.725 ;
        RECT 3.025 0.085 3.280 0.845 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__isobufsrc_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__isobufsrc_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__isobufsrc_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 4.845 1.075 5.425 1.320 ;
    END
  END A
  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.360 1.075 1.950 1.275 ;
    END
  END SLEEP
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.325 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.477000 ;
    PORT
      LAYER li1 ;
        RECT 2.545 1.745 2.715 2.125 ;
        RECT 3.485 1.745 3.655 2.125 ;
        RECT 2.545 1.445 3.655 1.745 ;
        RECT 2.545 0.905 2.875 1.445 ;
        RECT 0.535 0.725 3.735 0.905 ;
        RECT 0.535 0.255 0.915 0.725 ;
        RECT 1.475 0.255 1.855 0.725 ;
        RECT 2.415 0.255 2.795 0.725 ;
        RECT 3.355 0.255 3.735 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.085 1.665 0.365 2.465 ;
        RECT 0.535 1.835 0.915 2.635 ;
        RECT 1.135 1.665 1.305 2.465 ;
        RECT 1.475 1.835 1.775 2.635 ;
        RECT 1.945 2.295 4.255 2.465 ;
        RECT 1.945 1.665 2.325 2.295 ;
        RECT 2.885 1.935 3.265 2.295 ;
        RECT 0.085 1.455 2.325 1.665 ;
        RECT 3.825 1.575 4.255 2.295 ;
        RECT 4.425 1.575 4.755 2.465 ;
        RECT 4.425 1.275 4.675 1.575 ;
        RECT 4.975 1.495 5.380 2.635 ;
        RECT 3.095 1.075 4.675 1.275 ;
        RECT 0.085 0.085 0.365 0.905 ;
        RECT 1.135 0.085 1.305 0.555 ;
        RECT 2.075 0.085 2.245 0.555 ;
        RECT 3.015 0.085 3.185 0.555 ;
        RECT 3.955 0.085 4.245 0.905 ;
        RECT 4.425 0.815 4.675 1.075 ;
        RECT 4.425 0.255 4.755 0.815 ;
        RECT 4.975 0.085 5.265 0.905 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__isobufsrc_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__isobufsrc_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__isobufsrc_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.660 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.065 0.505 1.285 ;
        RECT 0.085 0.255 0.315 1.065 ;
    END
  END A
  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.220000 ;
    PORT
      LAYER li1 ;
        RECT 5.790 1.075 8.880 1.275 ;
    END
  END SLEEP
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.660 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.245 0.105 9.645 1.015 ;
        RECT 0.245 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.850 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.660 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.889000 ;
    PORT
      LAYER li1 ;
        RECT 5.975 1.615 6.225 2.125 ;
        RECT 6.915 1.615 7.165 2.125 ;
        RECT 7.855 1.615 8.105 2.125 ;
        RECT 8.795 1.615 9.045 2.125 ;
        RECT 5.975 1.445 9.565 1.615 ;
        RECT 9.050 0.905 9.565 1.445 ;
        RECT 2.125 0.725 9.565 0.905 ;
        RECT 2.125 0.255 2.505 0.725 ;
        RECT 3.065 0.255 3.445 0.725 ;
        RECT 4.005 0.255 4.385 0.725 ;
        RECT 4.945 0.255 5.325 0.725 ;
        RECT 5.885 0.255 6.265 0.725 ;
        RECT 6.825 0.255 7.205 0.725 ;
        RECT 7.765 0.255 8.145 0.725 ;
        RECT 8.705 0.255 9.085 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.660 2.805 ;
        RECT 0.125 1.455 0.345 2.635 ;
        RECT 0.515 1.455 0.945 2.465 ;
        RECT 1.165 1.455 1.460 2.635 ;
        RECT 1.675 1.665 1.995 2.465 ;
        RECT 2.215 1.835 2.465 2.635 ;
        RECT 2.685 1.665 2.935 2.465 ;
        RECT 3.155 1.835 3.405 2.635 ;
        RECT 3.625 1.665 3.875 2.465 ;
        RECT 4.095 1.835 4.345 2.635 ;
        RECT 4.565 1.665 4.815 2.465 ;
        RECT 5.035 1.835 5.285 2.635 ;
        RECT 5.505 2.295 9.515 2.465 ;
        RECT 5.505 1.665 5.755 2.295 ;
        RECT 6.445 1.785 6.695 2.295 ;
        RECT 7.385 1.785 7.635 2.295 ;
        RECT 8.325 1.785 8.575 2.295 ;
        RECT 9.265 1.785 9.515 2.295 ;
        RECT 1.675 1.455 5.755 1.665 ;
        RECT 0.725 1.285 0.945 1.455 ;
        RECT 0.725 1.075 5.520 1.285 ;
        RECT 0.725 1.065 1.235 1.075 ;
        RECT 0.485 0.085 0.705 0.895 ;
        RECT 0.875 0.255 1.235 1.065 ;
        RECT 1.445 0.085 1.955 0.905 ;
        RECT 2.725 0.085 2.895 0.555 ;
        RECT 3.665 0.085 3.835 0.555 ;
        RECT 4.605 0.085 4.775 0.555 ;
        RECT 5.545 0.085 5.715 0.555 ;
        RECT 6.485 0.085 6.655 0.555 ;
        RECT 7.425 0.085 7.595 0.555 ;
        RECT 8.365 0.085 8.535 0.555 ;
        RECT 9.305 0.085 9.575 0.555 ;
        RECT 0.000 -0.085 9.660 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__isobufsrc_8

#--------EOF---------

MACRO sky130_fd_sc_hdll__isobufsrc_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__isobufsrc_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.400 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.665 1.325 ;
        RECT 0.085 0.255 0.315 0.995 ;
    END
  END A
  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.440000 ;
    PORT
      LAYER li1 ;
        RECT 10.650 1.075 17.600 1.285 ;
    END
  END SLEEP
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 18.400 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 18.590 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 18.400 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.713000 ;
    PORT
      LAYER li1 ;
        RECT 10.935 1.625 11.185 2.125 ;
        RECT 11.875 1.625 12.125 2.125 ;
        RECT 12.815 1.625 13.065 2.125 ;
        RECT 13.755 1.625 14.005 2.125 ;
        RECT 14.695 1.625 14.945 2.125 ;
        RECT 15.635 1.625 15.885 2.125 ;
        RECT 16.575 1.625 16.825 2.125 ;
        RECT 17.515 1.625 17.765 2.125 ;
        RECT 10.935 1.455 18.305 1.625 ;
        RECT 17.770 0.905 18.305 1.455 ;
        RECT 3.325 0.725 18.305 0.905 ;
        RECT 3.325 0.255 3.705 0.725 ;
        RECT 4.265 0.255 4.645 0.725 ;
        RECT 5.205 0.255 5.585 0.725 ;
        RECT 6.145 0.255 6.525 0.725 ;
        RECT 7.085 0.255 7.465 0.725 ;
        RECT 8.025 0.255 8.405 0.725 ;
        RECT 8.965 0.255 9.345 0.725 ;
        RECT 9.905 0.255 10.285 0.725 ;
        RECT 10.845 0.255 11.225 0.725 ;
        RECT 11.785 0.255 12.165 0.725 ;
        RECT 12.725 0.255 13.105 0.725 ;
        RECT 13.665 0.255 14.045 0.725 ;
        RECT 14.605 0.255 14.985 0.725 ;
        RECT 15.545 0.255 15.925 0.725 ;
        RECT 16.485 0.255 16.865 0.725 ;
        RECT 17.425 0.255 17.805 0.725 ;
    END
  END X
  OBS
      LAYER pwell ;
        RECT 0.395 0.105 18.365 1.015 ;
      LAYER li1 ;
        RECT 0.000 2.635 18.400 2.805 ;
        RECT 0.300 1.495 0.515 2.635 ;
        RECT 0.685 1.495 1.115 2.465 ;
        RECT 0.885 1.285 1.115 1.495 ;
        RECT 1.335 1.455 1.555 2.635 ;
        RECT 1.725 1.285 2.155 2.465 ;
        RECT 2.375 1.455 2.670 2.635 ;
        RECT 2.875 1.665 3.195 2.465 ;
        RECT 3.415 1.835 3.665 2.635 ;
        RECT 3.885 1.665 4.135 2.465 ;
        RECT 4.355 1.835 4.605 2.635 ;
        RECT 4.825 1.665 5.075 2.465 ;
        RECT 5.295 1.835 5.545 2.635 ;
        RECT 5.765 1.665 6.015 2.465 ;
        RECT 6.235 1.835 6.485 2.635 ;
        RECT 6.705 1.665 6.955 2.465 ;
        RECT 7.175 1.835 7.425 2.635 ;
        RECT 7.645 1.665 7.895 2.465 ;
        RECT 8.115 1.835 8.365 2.635 ;
        RECT 8.585 1.665 8.835 2.465 ;
        RECT 9.055 1.835 9.305 2.635 ;
        RECT 9.525 1.665 9.775 2.465 ;
        RECT 9.995 1.835 10.245 2.635 ;
        RECT 10.465 2.295 18.235 2.465 ;
        RECT 10.465 1.665 10.715 2.295 ;
        RECT 11.405 1.795 11.655 2.295 ;
        RECT 12.345 1.795 12.595 2.295 ;
        RECT 13.285 1.795 13.535 2.295 ;
        RECT 14.225 1.795 14.475 2.295 ;
        RECT 15.165 1.795 15.415 2.295 ;
        RECT 16.105 1.795 16.355 2.295 ;
        RECT 17.045 1.795 17.295 2.295 ;
        RECT 17.985 1.795 18.235 2.295 ;
        RECT 2.875 1.455 10.715 1.665 ;
        RECT 0.885 1.075 10.480 1.285 ;
        RECT 0.885 1.065 2.385 1.075 ;
        RECT 0.485 0.085 0.865 0.825 ;
        RECT 1.085 0.255 1.345 1.065 ;
        RECT 1.565 0.085 1.865 0.895 ;
        RECT 2.085 0.255 2.385 1.065 ;
        RECT 2.605 0.085 3.155 0.905 ;
        RECT 3.925 0.085 4.095 0.555 ;
        RECT 4.865 0.085 5.035 0.555 ;
        RECT 5.805 0.085 5.975 0.555 ;
        RECT 6.745 0.085 6.915 0.555 ;
        RECT 7.685 0.085 7.855 0.555 ;
        RECT 8.625 0.085 8.795 0.555 ;
        RECT 9.565 0.085 9.735 0.555 ;
        RECT 10.505 0.085 10.675 0.555 ;
        RECT 11.445 0.085 11.615 0.555 ;
        RECT 12.385 0.085 12.555 0.555 ;
        RECT 13.325 0.085 13.495 0.555 ;
        RECT 14.265 0.085 14.435 0.555 ;
        RECT 15.205 0.085 15.375 0.555 ;
        RECT 16.145 0.085 16.315 0.555 ;
        RECT 17.085 0.085 17.255 0.555 ;
        RECT 18.025 0.085 18.295 0.555 ;
        RECT 0.000 -0.085 18.400 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 14.405 2.635 14.575 2.805 ;
        RECT 14.865 2.635 15.035 2.805 ;
        RECT 15.325 2.635 15.495 2.805 ;
        RECT 15.785 2.635 15.955 2.805 ;
        RECT 16.245 2.635 16.415 2.805 ;
        RECT 16.705 2.635 16.875 2.805 ;
        RECT 17.165 2.635 17.335 2.805 ;
        RECT 17.625 2.635 17.795 2.805 ;
        RECT 18.085 2.635 18.255 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
        RECT 14.405 -0.085 14.575 0.085 ;
        RECT 14.865 -0.085 15.035 0.085 ;
        RECT 15.325 -0.085 15.495 0.085 ;
        RECT 15.785 -0.085 15.955 0.085 ;
        RECT 16.245 -0.085 16.415 0.085 ;
        RECT 16.705 -0.085 16.875 0.085 ;
        RECT 17.165 -0.085 17.335 0.085 ;
        RECT 17.625 -0.085 17.795 0.085 ;
        RECT 18.085 -0.085 18.255 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__isobufsrc_16

#--------EOF---------

MACRO sky130_fd_sc_hdll__mux2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__mux2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 2.290 0.255 2.615 1.415 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.780 1.615 3.075 1.785 ;
        RECT 1.780 0.815 1.950 1.615 ;
        RECT 2.855 0.255 3.075 1.615 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277200 ;
    PORT
      LAYER li1 ;
        RECT 1.070 2.295 3.415 2.465 ;
        RECT 1.070 1.325 1.270 2.295 ;
        RECT 3.245 1.630 3.415 2.295 ;
        RECT 3.245 1.440 4.045 1.630 ;
        RECT 0.995 0.995 1.270 1.325 ;
    END
  END S
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.785 0.985 1.015 ;
        RECT 0.005 0.105 4.405 0.785 ;
        RECT 0.420 -0.085 0.640 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.495 0.425 2.465 ;
        RECT 0.090 0.255 0.345 1.495 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.645 1.495 0.815 2.635 ;
        RECT 1.440 1.955 2.750 2.125 ;
        RECT 0.515 0.825 0.685 1.325 ;
        RECT 1.440 0.825 1.610 1.955 ;
        RECT 3.585 1.875 3.755 2.635 ;
        RECT 4.040 1.875 4.500 2.285 ;
        RECT 4.215 1.065 4.500 1.875 ;
        RECT 3.285 0.895 4.500 1.065 ;
        RECT 0.515 0.655 1.610 0.825 ;
        RECT 1.435 0.620 1.610 0.655 ;
        RECT 0.515 0.085 0.895 0.485 ;
        RECT 1.435 0.255 1.955 0.620 ;
        RECT 3.250 0.085 3.765 0.620 ;
        RECT 4.035 0.290 4.280 0.895 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__mux2_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__mux2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__mux2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 2.135 1.410 3.075 1.625 ;
        RECT 2.125 1.325 3.075 1.410 ;
        RECT 1.920 1.280 3.075 1.325 ;
        RECT 1.920 0.765 2.295 1.280 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 2.530 0.775 3.075 1.105 ;
        RECT 2.870 0.420 3.075 0.775 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.356400 ;
    PORT
      LAYER li1 ;
        RECT 3.355 0.755 3.545 1.625 ;
    END
  END S
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.785 1.445 1.015 ;
        RECT 0.005 0.105 4.325 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.498000 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.595 0.875 2.465 ;
        RECT 0.515 0.255 0.800 1.595 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.090 1.495 0.345 2.635 ;
        RECT 1.115 2.175 1.285 2.635 ;
        RECT 1.455 2.255 2.860 2.425 ;
        RECT 1.455 2.005 1.625 2.255 ;
        RECT 3.460 2.175 3.680 2.635 ;
        RECT 3.850 2.005 4.235 2.465 ;
        RECT 1.095 1.835 1.625 2.005 ;
        RECT 1.795 1.835 4.235 2.005 ;
        RECT 1.095 1.325 1.265 1.835 ;
        RECT 1.795 1.665 1.965 1.835 ;
        RECT 0.970 0.995 1.265 1.325 ;
        RECT 1.435 1.495 1.965 1.665 ;
        RECT 1.435 0.995 1.655 1.495 ;
        RECT 0.090 0.085 0.345 0.885 ;
        RECT 1.095 0.805 1.265 0.995 ;
        RECT 1.095 0.635 1.705 0.805 ;
        RECT 1.535 0.595 1.705 0.635 ;
        RECT 0.985 0.085 1.365 0.465 ;
        RECT 1.535 0.265 2.250 0.595 ;
        RECT 3.485 0.085 3.685 0.585 ;
        RECT 3.985 0.255 4.235 1.835 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__mux2_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__mux2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__mux2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.450 0.995 1.795 1.615 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.965 0.995 2.585 1.325 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.430 0.995 0.790 1.325 ;
        RECT 0.620 0.805 0.790 0.995 ;
        RECT 2.880 0.995 3.595 1.325 ;
        RECT 2.880 0.805 3.050 0.995 ;
        RECT 0.620 0.635 3.050 0.805 ;
    END
  END S
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.965 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.996000 ;
    PORT
      LAYER li1 ;
        RECT 4.215 1.745 4.385 2.465 ;
        RECT 5.155 1.745 5.325 2.465 ;
        RECT 4.215 1.575 5.880 1.745 ;
        RECT 5.650 0.805 5.880 1.575 ;
        RECT 4.215 0.635 5.880 0.805 ;
        RECT 4.215 0.255 4.385 0.635 ;
        RECT 5.155 0.255 5.325 0.635 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.090 1.665 0.345 2.465 ;
        RECT 0.515 1.835 0.870 2.635 ;
        RECT 1.040 2.275 2.970 2.445 ;
        RECT 1.040 1.935 1.440 2.275 ;
        RECT 3.275 2.105 3.445 2.465 ;
        RECT 3.615 2.255 3.995 2.635 ;
        RECT 1.630 1.935 3.445 2.105 ;
        RECT 4.555 1.915 4.935 2.635 ;
        RECT 5.495 1.915 5.875 2.635 ;
        RECT 0.090 1.495 1.180 1.665 ;
        RECT 2.130 1.595 3.985 1.765 ;
        RECT 0.090 0.625 0.260 1.495 ;
        RECT 0.960 0.995 1.180 1.495 ;
        RECT 3.815 1.245 3.985 1.595 ;
        RECT 3.815 1.075 5.430 1.245 ;
        RECT 3.815 0.825 3.985 1.075 ;
        RECT 3.260 0.655 3.985 0.825 ;
        RECT 0.090 0.295 0.345 0.625 ;
        RECT 3.260 0.465 3.430 0.655 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 2.075 0.295 3.430 0.465 ;
        RECT 3.615 0.085 3.995 0.465 ;
        RECT 4.555 0.085 4.935 0.465 ;
        RECT 5.495 0.085 5.875 0.465 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__mux2_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__mux2_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__mux2_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.580 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.552000 ;
    PORT
      LAYER li1 ;
        RECT 5.580 0.815 5.800 1.325 ;
        RECT 7.625 1.165 7.845 1.325 ;
        RECT 7.325 0.995 7.845 1.165 ;
        RECT 7.325 0.815 7.495 0.995 ;
        RECT 5.580 0.645 7.495 0.815 ;
        RECT 5.755 0.425 6.390 0.645 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.552000 ;
    PORT
      LAYER met1 ;
        RECT 4.620 1.260 4.960 1.305 ;
        RECT 8.765 1.260 9.115 1.305 ;
        RECT 4.620 1.120 9.115 1.260 ;
        RECT 4.620 1.075 4.960 1.120 ;
        RECT 8.765 1.075 9.115 1.120 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.829500 ;
    PORT
      LAYER met1 ;
        RECT 6.110 1.600 6.400 1.645 ;
        RECT 9.745 1.600 10.035 1.645 ;
        RECT 6.110 1.460 10.035 1.600 ;
        RECT 6.110 1.415 6.400 1.460 ;
        RECT 9.745 1.415 10.035 1.460 ;
    END
  END S
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.580 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.005 4.265 1.015 ;
        RECT 9.585 1.005 10.555 1.015 ;
        RECT 0.005 0.105 10.555 1.005 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.770 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.580 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.024500 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.745 0.815 2.465 ;
        RECT 1.585 1.745 1.755 2.465 ;
        RECT 2.525 1.745 2.695 2.465 ;
        RECT 3.465 1.745 3.635 2.465 ;
        RECT 0.605 1.575 3.635 1.745 ;
        RECT 0.605 0.805 0.865 1.575 ;
        RECT 0.605 0.635 3.635 0.805 ;
        RECT 0.605 0.255 0.815 0.635 ;
        RECT 1.585 0.295 1.755 0.635 ;
        RECT 2.525 0.255 2.695 0.635 ;
        RECT 3.465 0.295 3.635 0.635 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.580 2.805 ;
        RECT 0.090 1.915 0.425 2.635 ;
        RECT 0.985 1.915 1.365 2.635 ;
        RECT 1.925 1.915 2.305 2.635 ;
        RECT 2.865 1.915 3.245 2.635 ;
        RECT 3.805 2.255 4.185 2.635 ;
        RECT 4.630 2.255 6.405 2.425 ;
        RECT 6.675 2.175 6.845 2.635 ;
        RECT 7.030 2.255 9.445 2.425 ;
        RECT 9.665 2.255 10.045 2.635 ;
        RECT 10.215 2.085 10.385 2.465 ;
        RECT 3.805 1.835 8.975 2.005 ;
        RECT 9.415 1.915 10.385 2.085 ;
        RECT 3.805 1.245 3.975 1.835 ;
        RECT 9.415 1.665 9.635 1.915 ;
        RECT 10.215 1.795 10.385 1.915 ;
        RECT 1.085 1.075 3.975 1.245 ;
        RECT 3.805 0.805 3.975 1.075 ;
        RECT 4.145 1.495 6.585 1.665 ;
        RECT 4.145 0.995 4.365 1.495 ;
        RECT 4.705 1.275 4.925 1.325 ;
        RECT 4.690 1.105 4.925 1.275 ;
        RECT 4.705 0.995 4.925 1.105 ;
        RECT 6.170 0.995 6.585 1.495 ;
        RECT 6.895 1.495 9.635 1.665 ;
        RECT 6.895 0.995 7.115 1.495 ;
        RECT 8.885 0.995 9.170 1.325 ;
        RECT 5.170 0.805 5.340 0.935 ;
        RECT 8.150 0.805 8.370 0.935 ;
        RECT 3.805 0.635 5.340 0.805 ;
        RECT 7.715 0.635 8.370 0.805 ;
        RECT 9.415 0.815 9.635 1.495 ;
        RECT 9.805 0.995 10.235 1.615 ;
        RECT 9.415 0.645 10.385 0.815 ;
        RECT 0.090 0.085 0.425 0.465 ;
        RECT 0.985 0.085 1.365 0.465 ;
        RECT 1.925 0.085 2.305 0.465 ;
        RECT 2.865 0.085 3.245 0.465 ;
        RECT 3.805 0.085 4.185 0.465 ;
        RECT 4.355 0.295 5.525 0.465 ;
        RECT 6.660 0.085 6.990 0.465 ;
        RECT 7.175 0.295 8.565 0.465 ;
        RECT 9.665 0.085 10.045 0.465 ;
        RECT 10.215 0.295 10.385 0.645 ;
        RECT 0.000 -0.085 10.580 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 6.170 1.445 6.340 1.615 ;
        RECT 4.690 1.105 4.860 1.275 ;
        RECT 8.885 1.105 9.055 1.275 ;
        RECT 5.170 0.765 5.340 0.935 ;
        RECT 8.150 0.765 8.320 0.935 ;
        RECT 9.805 1.445 9.975 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
      LAYER met1 ;
        RECT 5.110 0.920 5.400 0.965 ;
        RECT 8.090 0.920 8.430 0.965 ;
        RECT 5.110 0.780 8.430 0.920 ;
        RECT 5.110 0.735 5.400 0.780 ;
        RECT 8.090 0.735 8.430 0.780 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__mux2_8

#--------EOF---------

MACRO sky130_fd_sc_hdll__mux2_12
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__mux2_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.560 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 8.105 1.075 9.455 1.325 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.565 1.075 1.915 1.325 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.665000 ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.075 4.275 1.325 ;
    END
  END S
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 16.560 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 16.175 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 16.750 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 16.560 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.793000 ;
    PORT
      LAYER li1 ;
        RECT 10.585 1.665 10.915 2.465 ;
        RECT 11.525 1.665 11.855 2.465 ;
        RECT 12.465 1.665 12.795 2.465 ;
        RECT 13.405 1.665 13.735 2.465 ;
        RECT 14.345 1.665 14.675 2.465 ;
        RECT 15.285 1.665 15.615 2.465 ;
        RECT 10.585 1.495 15.615 1.665 ;
        RECT 15.285 0.905 15.615 1.495 ;
        RECT 10.585 0.725 15.615 0.905 ;
        RECT 10.585 0.255 10.915 0.725 ;
        RECT 11.525 0.255 11.855 0.725 ;
        RECT 12.465 0.255 12.795 0.725 ;
        RECT 13.405 0.255 13.735 0.725 ;
        RECT 14.345 0.255 14.675 0.725 ;
        RECT 15.285 0.255 15.615 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 16.560 2.805 ;
        RECT 0.095 2.295 2.305 2.465 ;
        RECT 0.095 0.425 0.395 2.295 ;
        RECT 0.565 1.665 0.895 2.125 ;
        RECT 1.065 1.835 1.335 2.295 ;
        RECT 1.505 1.665 1.835 2.125 ;
        RECT 0.565 1.495 1.835 1.665 ;
        RECT 2.005 1.495 2.305 2.295 ;
        RECT 2.525 1.495 2.795 2.635 ;
        RECT 2.965 1.665 3.295 2.465 ;
        RECT 3.465 1.835 3.735 2.635 ;
        RECT 3.905 1.665 4.235 2.465 ;
        RECT 2.965 1.495 4.235 1.665 ;
        RECT 4.405 1.495 4.675 2.635 ;
        RECT 4.845 1.325 5.175 2.465 ;
        RECT 5.345 1.495 5.615 2.635 ;
        RECT 5.785 1.665 6.115 2.465 ;
        RECT 6.285 1.835 6.555 2.635 ;
        RECT 6.725 1.665 7.055 2.465 ;
        RECT 5.785 1.495 7.055 1.665 ;
        RECT 7.225 1.495 7.495 2.635 ;
        RECT 7.715 2.295 9.925 2.465 ;
        RECT 7.715 1.495 8.015 2.295 ;
        RECT 8.185 1.665 8.515 2.125 ;
        RECT 8.685 1.835 8.955 2.295 ;
        RECT 9.125 1.665 9.455 2.125 ;
        RECT 8.185 1.495 9.455 1.665 ;
        RECT 9.625 1.325 9.925 2.295 ;
        RECT 10.145 1.495 10.415 2.635 ;
        RECT 11.085 1.835 11.355 2.635 ;
        RECT 12.025 1.835 12.295 2.635 ;
        RECT 12.965 1.835 13.235 2.635 ;
        RECT 13.905 1.835 14.175 2.635 ;
        RECT 14.845 1.835 15.115 2.635 ;
        RECT 15.785 1.495 16.055 2.635 ;
        RECT 4.845 1.075 7.095 1.325 ;
        RECT 9.625 1.075 14.825 1.325 ;
        RECT 0.565 0.725 4.235 0.905 ;
        RECT 0.565 0.595 0.895 0.725 ;
        RECT 1.505 0.595 1.835 0.725 ;
        RECT 1.065 0.425 1.335 0.545 ;
        RECT 2.005 0.425 2.305 0.550 ;
        RECT 0.095 0.255 2.305 0.425 ;
        RECT 2.525 0.085 2.795 0.550 ;
        RECT 2.965 0.255 3.295 0.725 ;
        RECT 3.465 0.085 3.735 0.545 ;
        RECT 3.905 0.255 4.235 0.725 ;
        RECT 4.405 0.085 4.675 0.905 ;
        RECT 4.845 0.255 5.175 1.075 ;
        RECT 5.345 0.085 5.615 0.905 ;
        RECT 5.785 0.725 9.455 0.905 ;
        RECT 5.785 0.255 6.115 0.725 ;
        RECT 6.285 0.085 6.555 0.545 ;
        RECT 6.725 0.255 7.055 0.725 ;
        RECT 8.185 0.595 8.515 0.725 ;
        RECT 9.125 0.595 9.455 0.725 ;
        RECT 7.225 0.085 7.495 0.550 ;
        RECT 7.715 0.425 8.015 0.550 ;
        RECT 8.685 0.425 8.955 0.545 ;
        RECT 9.625 0.425 9.925 1.075 ;
        RECT 7.715 0.255 9.925 0.425 ;
        RECT 10.145 0.085 10.415 0.905 ;
        RECT 11.085 0.085 11.355 0.545 ;
        RECT 12.025 0.085 12.295 0.545 ;
        RECT 12.965 0.085 13.235 0.545 ;
        RECT 13.905 0.085 14.175 0.550 ;
        RECT 14.845 0.085 15.115 0.545 ;
        RECT 15.785 0.085 16.055 0.905 ;
        RECT 0.000 -0.085 16.560 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 14.405 2.635 14.575 2.805 ;
        RECT 14.865 2.635 15.035 2.805 ;
        RECT 15.325 2.635 15.495 2.805 ;
        RECT 15.785 2.635 15.955 2.805 ;
        RECT 16.245 2.635 16.415 2.805 ;
        RECT 0.645 1.785 0.815 1.955 ;
        RECT 1.585 1.785 1.755 1.955 ;
        RECT 3.045 2.125 3.215 2.295 ;
        RECT 3.985 2.125 4.155 2.295 ;
        RECT 5.865 1.785 6.035 1.955 ;
        RECT 6.805 1.785 6.975 1.955 ;
        RECT 8.265 1.785 8.435 1.955 ;
        RECT 9.205 1.785 9.375 1.955 ;
        RECT 0.175 0.425 0.345 0.595 ;
        RECT 9.675 0.425 9.845 0.595 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
        RECT 14.405 -0.085 14.575 0.085 ;
        RECT 14.865 -0.085 15.035 0.085 ;
        RECT 15.325 -0.085 15.495 0.085 ;
        RECT 15.785 -0.085 15.955 0.085 ;
        RECT 16.245 -0.085 16.415 0.085 ;
      LAYER met1 ;
        RECT 2.985 2.280 3.275 2.325 ;
        RECT 3.925 2.280 4.215 2.325 ;
        RECT 2.985 2.140 7.660 2.280 ;
        RECT 2.985 2.095 3.275 2.140 ;
        RECT 3.925 2.095 4.215 2.140 ;
        RECT 0.585 1.940 0.875 1.985 ;
        RECT 1.525 1.940 1.815 1.985 ;
        RECT 5.805 1.940 6.095 1.985 ;
        RECT 6.745 1.940 7.035 1.985 ;
        RECT 0.585 1.800 7.035 1.940 ;
        RECT 7.520 1.940 7.660 2.140 ;
        RECT 8.205 1.940 8.495 1.985 ;
        RECT 9.145 1.940 9.435 1.985 ;
        RECT 7.520 1.800 9.435 1.940 ;
        RECT 0.585 1.755 0.875 1.800 ;
        RECT 1.525 1.755 1.815 1.800 ;
        RECT 5.805 1.755 6.095 1.800 ;
        RECT 6.745 1.755 7.035 1.800 ;
        RECT 8.205 1.755 8.495 1.800 ;
        RECT 9.145 1.755 9.435 1.800 ;
        RECT 0.115 0.580 0.405 0.625 ;
        RECT 9.615 0.580 9.905 0.625 ;
        RECT 0.115 0.440 9.905 0.580 ;
        RECT 0.115 0.395 0.405 0.440 ;
        RECT 9.615 0.395 9.905 0.440 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__mux2_12

#--------EOF---------

MACRO sky130_fd_sc_hdll__mux2_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__mux2_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.400 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 8.105 1.075 9.455 1.325 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.565 1.075 1.915 1.325 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.665000 ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.075 4.275 1.325 ;
    END
  END S
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 18.400 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 18.055 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 18.590 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 18.400 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.724000 ;
    PORT
      LAYER li1 ;
        RECT 10.585 1.665 10.915 2.465 ;
        RECT 11.525 1.665 11.855 2.465 ;
        RECT 12.465 1.665 12.795 2.465 ;
        RECT 13.405 1.665 13.735 2.465 ;
        RECT 14.345 1.665 14.675 2.465 ;
        RECT 15.285 1.665 15.615 2.465 ;
        RECT 16.225 1.665 16.555 2.465 ;
        RECT 17.165 1.665 17.495 2.465 ;
        RECT 10.585 1.495 17.495 1.665 ;
        RECT 17.085 0.905 17.495 1.495 ;
        RECT 10.585 0.725 17.495 0.905 ;
        RECT 10.585 0.255 10.915 0.725 ;
        RECT 11.525 0.255 11.855 0.725 ;
        RECT 12.465 0.255 12.795 0.725 ;
        RECT 13.405 0.255 13.735 0.725 ;
        RECT 14.345 0.255 14.675 0.725 ;
        RECT 15.285 0.255 15.615 0.725 ;
        RECT 16.225 0.255 16.555 0.725 ;
        RECT 17.165 0.255 17.495 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 18.400 2.805 ;
        RECT 0.095 2.295 2.305 2.465 ;
        RECT 0.095 0.425 0.395 2.295 ;
        RECT 0.565 1.665 0.895 2.125 ;
        RECT 1.065 1.835 1.335 2.295 ;
        RECT 1.505 1.665 1.835 2.125 ;
        RECT 0.565 1.495 1.835 1.665 ;
        RECT 2.005 1.495 2.305 2.295 ;
        RECT 2.525 1.495 2.795 2.635 ;
        RECT 2.965 1.665 3.295 2.465 ;
        RECT 3.465 1.835 3.735 2.635 ;
        RECT 3.905 1.665 4.235 2.465 ;
        RECT 2.965 1.495 4.235 1.665 ;
        RECT 4.405 1.495 4.675 2.635 ;
        RECT 4.845 1.325 5.175 2.465 ;
        RECT 5.345 1.495 5.615 2.635 ;
        RECT 5.785 1.665 6.115 2.465 ;
        RECT 6.285 1.835 6.555 2.635 ;
        RECT 6.725 1.665 7.055 2.465 ;
        RECT 5.785 1.495 7.055 1.665 ;
        RECT 7.225 1.495 7.495 2.635 ;
        RECT 7.715 2.295 9.925 2.465 ;
        RECT 7.715 1.495 8.015 2.295 ;
        RECT 8.185 1.665 8.515 2.125 ;
        RECT 8.685 1.835 8.955 2.295 ;
        RECT 9.125 1.665 9.455 2.125 ;
        RECT 8.185 1.495 9.455 1.665 ;
        RECT 9.625 1.325 9.925 2.295 ;
        RECT 10.145 1.495 10.415 2.635 ;
        RECT 11.085 1.835 11.355 2.635 ;
        RECT 12.025 1.835 12.295 2.635 ;
        RECT 12.965 1.835 13.235 2.635 ;
        RECT 13.905 1.835 14.175 2.635 ;
        RECT 14.845 1.835 15.115 2.635 ;
        RECT 15.785 1.835 16.055 2.635 ;
        RECT 16.725 1.835 16.995 2.635 ;
        RECT 17.665 1.495 17.935 2.635 ;
        RECT 4.845 1.075 7.095 1.325 ;
        RECT 9.625 1.075 16.865 1.325 ;
        RECT 0.565 0.725 4.235 0.905 ;
        RECT 0.565 0.595 0.895 0.725 ;
        RECT 1.505 0.595 1.835 0.725 ;
        RECT 1.065 0.425 1.335 0.545 ;
        RECT 2.005 0.425 2.305 0.550 ;
        RECT 0.095 0.255 2.305 0.425 ;
        RECT 2.525 0.085 2.795 0.550 ;
        RECT 2.965 0.255 3.295 0.725 ;
        RECT 3.465 0.085 3.735 0.545 ;
        RECT 3.905 0.255 4.235 0.725 ;
        RECT 4.405 0.085 4.675 0.905 ;
        RECT 4.845 0.255 5.175 1.075 ;
        RECT 5.345 0.085 5.615 0.905 ;
        RECT 5.785 0.725 9.455 0.905 ;
        RECT 5.785 0.255 6.115 0.725 ;
        RECT 6.285 0.085 6.555 0.545 ;
        RECT 6.725 0.255 7.055 0.725 ;
        RECT 8.185 0.595 8.515 0.725 ;
        RECT 9.125 0.595 9.455 0.725 ;
        RECT 7.225 0.085 7.495 0.550 ;
        RECT 7.715 0.425 8.015 0.550 ;
        RECT 8.685 0.425 8.955 0.545 ;
        RECT 9.625 0.425 9.925 1.075 ;
        RECT 7.715 0.255 9.925 0.425 ;
        RECT 10.145 0.085 10.415 0.905 ;
        RECT 11.085 0.085 11.355 0.545 ;
        RECT 12.025 0.085 12.295 0.545 ;
        RECT 12.965 0.085 13.235 0.545 ;
        RECT 13.905 0.085 14.175 0.550 ;
        RECT 14.845 0.085 15.115 0.545 ;
        RECT 15.785 0.085 16.055 0.545 ;
        RECT 16.725 0.085 16.995 0.545 ;
        RECT 17.665 0.085 17.935 0.905 ;
        RECT 0.000 -0.085 18.400 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 14.405 2.635 14.575 2.805 ;
        RECT 14.865 2.635 15.035 2.805 ;
        RECT 15.325 2.635 15.495 2.805 ;
        RECT 15.785 2.635 15.955 2.805 ;
        RECT 16.245 2.635 16.415 2.805 ;
        RECT 16.705 2.635 16.875 2.805 ;
        RECT 17.165 2.635 17.335 2.805 ;
        RECT 17.625 2.635 17.795 2.805 ;
        RECT 18.085 2.635 18.255 2.805 ;
        RECT 0.645 1.785 0.815 1.955 ;
        RECT 1.585 1.785 1.755 1.955 ;
        RECT 3.045 2.125 3.215 2.295 ;
        RECT 3.985 2.125 4.155 2.295 ;
        RECT 5.865 1.785 6.035 1.955 ;
        RECT 6.805 1.785 6.975 1.955 ;
        RECT 8.265 1.785 8.435 1.955 ;
        RECT 9.205 1.785 9.375 1.955 ;
        RECT 0.175 0.425 0.345 0.595 ;
        RECT 9.675 0.425 9.845 0.595 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
        RECT 14.405 -0.085 14.575 0.085 ;
        RECT 14.865 -0.085 15.035 0.085 ;
        RECT 15.325 -0.085 15.495 0.085 ;
        RECT 15.785 -0.085 15.955 0.085 ;
        RECT 16.245 -0.085 16.415 0.085 ;
        RECT 16.705 -0.085 16.875 0.085 ;
        RECT 17.165 -0.085 17.335 0.085 ;
        RECT 17.625 -0.085 17.795 0.085 ;
        RECT 18.085 -0.085 18.255 0.085 ;
      LAYER met1 ;
        RECT 2.985 2.280 3.275 2.325 ;
        RECT 3.925 2.280 4.215 2.325 ;
        RECT 2.985 2.140 7.660 2.280 ;
        RECT 2.985 2.095 3.275 2.140 ;
        RECT 3.925 2.095 4.215 2.140 ;
        RECT 0.585 1.940 0.875 1.985 ;
        RECT 1.525 1.940 1.815 1.985 ;
        RECT 5.805 1.940 6.095 1.985 ;
        RECT 6.745 1.940 7.035 1.985 ;
        RECT 0.585 1.800 7.035 1.940 ;
        RECT 7.520 1.940 7.660 2.140 ;
        RECT 8.205 1.940 8.495 1.985 ;
        RECT 9.145 1.940 9.435 1.985 ;
        RECT 7.520 1.800 9.435 1.940 ;
        RECT 0.585 1.755 0.875 1.800 ;
        RECT 1.525 1.755 1.815 1.800 ;
        RECT 5.805 1.755 6.095 1.800 ;
        RECT 6.745 1.755 7.035 1.800 ;
        RECT 8.205 1.755 8.495 1.800 ;
        RECT 9.145 1.755 9.435 1.800 ;
        RECT 0.115 0.580 0.405 0.625 ;
        RECT 9.615 0.580 9.905 0.625 ;
        RECT 0.115 0.440 9.905 0.580 ;
        RECT 0.115 0.395 0.405 0.440 ;
        RECT 9.615 0.395 9.905 0.440 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__mux2_16

#--------EOF---------

MACRO sky130_fd_sc_hdll__mux2i_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__mux2i_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.060 0.420 1.285 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.325 1.265 2.110 ;
        RECT 1.005 0.995 1.265 1.325 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 3.365 0.760 3.750 1.620 ;
    END
  END S
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.855 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.465500 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.455 0.890 2.125 ;
        RECT 0.605 0.595 0.835 1.455 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.120 2.295 1.725 2.465 ;
        RECT 0.120 1.455 0.420 2.295 ;
        RECT 1.505 1.650 1.725 2.295 ;
        RECT 1.895 1.835 2.175 2.635 ;
        RECT 2.365 1.650 2.745 2.465 ;
        RECT 1.505 1.480 2.745 1.650 ;
        RECT 2.970 1.310 3.195 2.465 ;
        RECT 3.475 1.835 3.770 2.635 ;
        RECT 1.485 1.075 3.195 1.310 ;
        RECT 0.085 0.465 0.345 0.885 ;
        RECT 1.575 0.825 2.700 0.885 ;
        RECT 1.005 0.715 2.700 0.825 ;
        RECT 1.005 0.655 1.750 0.715 ;
        RECT 0.085 0.425 0.440 0.465 ;
        RECT 1.065 0.425 1.855 0.465 ;
        RECT 0.085 0.255 1.855 0.425 ;
        RECT 2.025 0.085 2.195 0.525 ;
        RECT 2.465 0.255 2.700 0.715 ;
        RECT 2.930 0.255 3.195 1.075 ;
        RECT 3.515 0.085 3.735 0.545 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__mux2i_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__mux2i_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__mux2i_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.720 1.075 4.025 1.275 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 4.710 0.995 5.085 1.615 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.832500 ;
    PORT
      LAYER li1 ;
        RECT 0.430 0.995 0.830 1.325 ;
        RECT 0.630 0.725 0.830 0.995 ;
    END
  END S
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.505 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.796250 ;
    PORT
      LAYER li1 ;
        RECT 2.965 2.255 5.425 2.425 ;
        RECT 5.200 1.785 5.425 2.255 ;
        RECT 5.255 0.465 5.425 1.785 ;
        RECT 2.965 0.295 5.425 0.465 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.085 2.135 0.345 2.465 ;
        RECT 0.515 2.255 0.895 2.635 ;
        RECT 1.455 2.255 1.835 2.635 ;
        RECT 2.055 2.135 2.280 2.465 ;
        RECT 2.525 2.175 2.775 2.635 ;
        RECT 0.085 1.665 0.260 2.135 ;
        RECT 2.110 2.005 2.280 2.135 ;
        RECT 2.965 2.005 4.750 2.085 ;
        RECT 0.985 1.835 1.885 2.005 ;
        RECT 2.110 1.915 4.750 2.005 ;
        RECT 2.110 1.835 3.135 1.915 ;
        RECT 1.715 1.665 1.885 1.835 ;
        RECT 3.385 1.665 3.765 1.715 ;
        RECT 0.085 1.495 1.545 1.665 ;
        RECT 1.715 1.495 3.765 1.665 ;
        RECT 0.085 0.675 0.260 1.495 ;
        RECT 1.325 1.325 1.545 1.495 ;
        RECT 1.325 1.155 2.185 1.325 ;
        RECT 1.805 1.075 2.185 1.155 ;
        RECT 0.085 0.345 0.345 0.675 ;
        RECT 1.115 0.575 1.355 0.935 ;
        RECT 0.515 0.085 0.885 0.545 ;
        RECT 1.585 0.085 1.835 0.885 ;
        RECT 2.055 0.735 3.765 0.905 ;
        RECT 2.055 0.295 2.225 0.735 ;
        RECT 3.385 0.655 3.765 0.735 ;
        RECT 4.200 0.825 4.505 0.935 ;
        RECT 4.200 0.655 4.745 0.825 ;
        RECT 2.525 0.085 2.695 0.545 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 1.170 0.765 1.340 0.935 ;
        RECT 4.200 0.765 4.370 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
      LAYER met1 ;
        RECT 1.110 0.920 1.400 0.965 ;
        RECT 4.140 0.920 4.480 0.965 ;
        RECT 1.110 0.780 4.480 0.920 ;
        RECT 1.110 0.735 1.400 0.780 ;
        RECT 4.140 0.735 4.480 0.780 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__mux2i_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__mux2i_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__mux2i_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.200 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 0.995 1.235 1.325 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 2.355 0.995 4.050 1.325 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.387500 ;
    PORT
      LAYER li1 ;
        RECT 6.360 1.425 8.650 1.595 ;
        RECT 6.360 1.290 6.530 1.425 ;
        RECT 4.245 1.075 6.530 1.290 ;
        RECT 8.480 0.995 8.650 1.425 ;
    END
  END S
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.200 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 9.125 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.390 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.200 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.339500 ;
    PORT
      LAYER li1 ;
        RECT 0.095 2.255 4.185 2.425 ;
        RECT 0.095 0.485 0.320 2.255 ;
        RECT 0.095 0.315 4.185 0.485 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.200 2.805 ;
        RECT 4.375 2.255 4.705 2.635 ;
        RECT 5.265 2.255 5.645 2.635 ;
        RECT 6.205 2.255 6.585 2.635 ;
        RECT 6.805 2.085 6.975 2.465 ;
        RECT 7.145 2.255 7.525 2.635 ;
        RECT 7.745 2.085 7.915 2.465 ;
        RECT 8.235 2.255 8.565 2.635 ;
        RECT 2.395 1.915 7.915 2.085 ;
        RECT 6.805 1.795 6.975 1.915 ;
        RECT 7.745 1.795 7.915 1.915 ;
        RECT 8.785 1.795 9.045 2.465 ;
        RECT 0.515 1.575 6.130 1.745 ;
        RECT 7.430 1.075 8.310 1.245 ;
        RECT 1.455 0.825 1.850 0.935 ;
        RECT 6.800 0.905 7.100 0.935 ;
        RECT 0.515 0.655 1.850 0.825 ;
        RECT 2.395 0.655 6.035 0.825 ;
        RECT 4.375 0.085 4.705 0.465 ;
        RECT 4.925 0.255 5.095 0.655 ;
        RECT 5.265 0.085 5.645 0.465 ;
        RECT 5.865 0.255 6.035 0.655 ;
        RECT 6.800 0.715 7.915 0.905 ;
        RECT 6.205 0.085 6.580 0.590 ;
        RECT 6.800 0.255 6.975 0.715 ;
        RECT 7.245 0.085 7.495 0.545 ;
        RECT 7.745 0.510 7.915 0.715 ;
        RECT 8.090 0.825 8.310 1.075 ;
        RECT 8.870 0.825 9.045 1.795 ;
        RECT 8.090 0.655 9.045 0.825 ;
        RECT 8.235 0.085 8.565 0.465 ;
        RECT 8.785 0.255 9.045 0.655 ;
        RECT 0.000 -0.085 9.200 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 1.680 0.765 1.850 0.935 ;
        RECT 6.800 0.765 6.970 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
      LAYER met1 ;
        RECT 1.620 0.920 1.910 0.965 ;
        RECT 6.690 0.920 7.030 0.965 ;
        RECT 1.620 0.780 7.030 0.920 ;
        RECT 1.620 0.735 1.910 0.780 ;
        RECT 6.690 0.735 7.030 0.780 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__mux2i_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__muxb4to1_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__muxb4to1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.740 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 8.010 1.055 8.405 1.325 ;
        RECT 8.010 0.625 8.180 1.055 ;
        RECT 7.905 0.395 8.180 0.625 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 4.475 1.055 4.870 1.325 ;
        RECT 4.700 0.625 4.870 1.055 ;
        RECT 4.700 0.395 4.975 0.625 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 3.870 1.055 4.265 1.325 ;
        RECT 3.870 0.625 4.040 1.055 ;
        RECT 3.765 0.395 4.040 0.625 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.335 1.055 0.730 1.325 ;
        RECT 0.560 0.625 0.730 1.055 ;
        RECT 0.560 0.395 0.835 0.625 ;
    END
  END D[0]
  PIN S[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 6.585 0.945 6.935 1.295 ;
    END
  END S[3]
  PIN S[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 5.945 0.945 6.295 1.295 ;
    END
  END S[2]
  PIN S[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 2.445 0.945 2.795 1.295 ;
    END
  END S[1]
  PIN S[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 1.805 0.945 2.155 1.295 ;
    END
  END S[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.740 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.885 0.925 1.015 ;
        RECT 3.675 0.885 5.065 1.015 ;
        RECT 7.815 0.885 8.735 1.015 ;
        RECT 0.005 0.105 8.735 0.885 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.930 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.740 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.426400 ;
    PORT
      LAYER met1 ;
        RECT 1.005 1.940 1.295 1.985 ;
        RECT 3.305 1.940 3.595 1.985 ;
        RECT 5.145 1.940 5.435 1.985 ;
        RECT 7.445 1.940 7.735 1.985 ;
        RECT 1.005 1.800 7.735 1.940 ;
        RECT 1.005 1.755 1.295 1.800 ;
        RECT 3.305 1.755 3.595 1.800 ;
        RECT 5.145 1.755 5.435 1.800 ;
        RECT 7.445 1.755 7.735 1.800 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.740 2.805 ;
        RECT 0.095 1.495 0.425 2.635 ;
        RECT 1.090 1.985 1.420 2.465 ;
        RECT 0.900 1.805 1.420 1.985 ;
        RECT 0.900 1.755 1.295 1.805 ;
        RECT 0.900 1.005 1.070 1.755 ;
        RECT 1.610 1.635 1.940 2.465 ;
        RECT 1.460 1.505 1.940 1.635 ;
        RECT 1.240 1.465 1.940 1.505 ;
        RECT 2.165 1.465 2.465 2.635 ;
        RECT 2.660 1.635 2.990 2.465 ;
        RECT 3.180 1.985 3.510 2.465 ;
        RECT 3.180 1.805 3.700 1.985 ;
        RECT 3.305 1.755 3.700 1.805 ;
        RECT 2.660 1.505 3.140 1.635 ;
        RECT 2.660 1.465 3.360 1.505 ;
        RECT 1.240 1.175 1.630 1.465 ;
        RECT 0.130 0.085 0.390 0.885 ;
        RECT 0.900 0.835 1.290 1.005 ;
        RECT 1.045 0.330 1.290 0.835 ;
        RECT 1.460 0.755 1.630 1.175 ;
        RECT 2.970 1.175 3.360 1.465 ;
        RECT 2.970 0.755 3.140 1.175 ;
        RECT 3.530 1.005 3.700 1.755 ;
        RECT 4.175 1.495 4.565 2.635 ;
        RECT 5.230 1.985 5.560 2.465 ;
        RECT 5.040 1.805 5.560 1.985 ;
        RECT 5.040 1.755 5.435 1.805 ;
        RECT 1.460 0.585 1.900 0.755 ;
        RECT 1.650 0.330 1.900 0.585 ;
        RECT 2.135 0.085 2.465 0.660 ;
        RECT 2.700 0.585 3.140 0.755 ;
        RECT 3.310 0.835 3.700 1.005 ;
        RECT 5.040 1.005 5.210 1.755 ;
        RECT 5.750 1.635 6.080 2.465 ;
        RECT 5.600 1.505 6.080 1.635 ;
        RECT 5.380 1.465 6.080 1.505 ;
        RECT 6.275 1.465 6.575 2.635 ;
        RECT 6.800 1.635 7.130 2.465 ;
        RECT 7.320 1.985 7.650 2.465 ;
        RECT 7.320 1.805 7.840 1.985 ;
        RECT 7.445 1.755 7.840 1.805 ;
        RECT 6.800 1.505 7.280 1.635 ;
        RECT 6.800 1.465 7.500 1.505 ;
        RECT 5.380 1.175 5.770 1.465 ;
        RECT 2.700 0.330 2.950 0.585 ;
        RECT 3.310 0.330 3.555 0.835 ;
        RECT 4.210 0.085 4.530 0.885 ;
        RECT 5.040 0.835 5.430 1.005 ;
        RECT 5.185 0.330 5.430 0.835 ;
        RECT 5.600 0.755 5.770 1.175 ;
        RECT 7.110 1.175 7.500 1.465 ;
        RECT 7.110 0.755 7.280 1.175 ;
        RECT 7.670 1.005 7.840 1.755 ;
        RECT 8.315 1.495 8.645 2.635 ;
        RECT 5.600 0.585 6.040 0.755 ;
        RECT 5.790 0.330 6.040 0.585 ;
        RECT 6.275 0.085 6.605 0.660 ;
        RECT 6.840 0.585 7.280 0.755 ;
        RECT 7.450 0.835 7.840 1.005 ;
        RECT 6.840 0.330 7.090 0.585 ;
        RECT 7.450 0.330 7.695 0.835 ;
        RECT 8.350 0.085 8.610 0.885 ;
        RECT 0.000 -0.085 8.740 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 1.065 1.785 1.235 1.955 ;
        RECT 3.365 1.785 3.535 1.955 ;
        RECT 5.205 1.785 5.375 1.955 ;
        RECT 7.505 1.785 7.675 1.955 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__muxb4to1_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__muxb4to1_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__muxb4to1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.880 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 11.965 1.055 12.785 1.325 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 6.535 1.055 7.355 1.325 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 5.525 1.055 6.345 1.325 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.055 0.915 1.325 ;
    END
  END D[0]
  PIN S[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 9.755 1.025 10.090 1.295 ;
    END
  END S[3]
  PIN S[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 9.230 1.025 9.565 1.295 ;
    END
  END S[2]
  PIN S[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 3.315 1.025 3.650 1.295 ;
    END
  END S[1]
  PIN S[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 2.790 1.025 3.125 1.295 ;
    END
  END S[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 12.880 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.995 1.440 1.015 ;
        RECT 5.000 0.995 7.880 1.015 ;
        RECT 11.440 0.995 12.875 1.015 ;
        RECT 0.005 0.885 2.345 0.995 ;
        RECT 4.095 0.885 8.785 0.995 ;
        RECT 10.535 0.885 12.875 0.995 ;
        RECT 0.005 0.215 12.875 0.885 ;
        RECT 0.005 0.105 1.440 0.215 ;
        RECT 2.545 0.105 3.895 0.215 ;
        RECT 5.000 0.105 7.880 0.215 ;
        RECT 8.985 0.105 10.335 0.215 ;
        RECT 11.440 0.105 12.875 0.215 ;
        RECT 0.145 -0.085 0.315 0.105 ;
        RECT 6.125 -0.085 6.755 0.105 ;
        RECT 12.565 -0.085 12.735 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 13.070 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 12.880 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.512800 ;
    PORT
      LAYER met1 ;
        RECT 1.465 1.940 1.755 1.985 ;
        RECT 4.685 1.940 4.975 1.985 ;
        RECT 7.905 1.940 8.195 1.985 ;
        RECT 11.125 1.940 11.415 1.985 ;
        RECT 1.465 1.800 11.415 1.940 ;
        RECT 1.465 1.755 1.755 1.800 ;
        RECT 4.685 1.755 4.975 1.800 ;
        RECT 7.905 1.755 8.195 1.800 ;
        RECT 11.125 1.755 11.415 1.800 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 12.880 2.805 ;
        RECT 0.095 2.210 0.425 2.465 ;
        RECT 0.095 1.665 0.395 2.210 ;
        RECT 0.595 2.105 0.895 2.635 ;
        RECT 0.565 1.835 0.895 2.105 ;
        RECT 1.115 2.295 2.280 2.465 ;
        RECT 1.115 1.665 1.285 2.295 ;
        RECT 1.465 1.755 1.895 2.125 ;
        RECT 0.095 1.495 1.285 1.665 ;
        RECT 1.030 0.885 1.335 0.925 ;
        RECT 1.585 0.885 1.755 1.755 ;
        RECT 2.110 1.645 2.280 2.295 ;
        RECT 2.550 1.635 2.880 2.465 ;
        RECT 2.450 1.475 2.880 1.635 ;
        RECT 2.100 1.465 2.880 1.475 ;
        RECT 3.055 1.465 3.385 2.635 ;
        RECT 3.560 1.635 3.890 2.465 ;
        RECT 4.160 2.295 5.325 2.465 ;
        RECT 4.160 1.645 4.330 2.295 ;
        RECT 4.545 1.755 4.975 2.125 ;
        RECT 3.560 1.475 3.990 1.635 ;
        RECT 3.560 1.465 4.340 1.475 ;
        RECT 2.100 1.305 2.620 1.465 ;
        RECT 3.820 1.305 4.340 1.465 ;
        RECT 2.100 1.205 2.515 1.305 ;
        RECT 0.145 0.715 1.335 0.885 ;
        RECT 0.145 0.255 0.475 0.715 ;
        RECT 0.645 0.085 0.860 0.545 ;
        RECT 1.030 0.425 1.335 0.715 ;
        RECT 1.505 0.595 1.835 0.885 ;
        RECT 2.005 0.425 2.175 0.770 ;
        RECT 2.345 0.755 2.515 1.205 ;
        RECT 3.925 1.205 4.340 1.305 ;
        RECT 3.925 0.755 4.095 1.205 ;
        RECT 4.685 0.885 4.855 1.755 ;
        RECT 5.155 1.665 5.325 2.295 ;
        RECT 5.545 2.105 5.845 2.635 ;
        RECT 6.015 2.210 6.345 2.465 ;
        RECT 5.545 1.835 5.875 2.105 ;
        RECT 6.045 1.665 6.345 2.210 ;
        RECT 5.155 1.495 6.345 1.665 ;
        RECT 6.535 2.210 6.865 2.465 ;
        RECT 6.535 1.665 6.835 2.210 ;
        RECT 7.035 2.105 7.335 2.635 ;
        RECT 7.005 1.835 7.335 2.105 ;
        RECT 7.555 2.295 8.720 2.465 ;
        RECT 7.555 1.665 7.725 2.295 ;
        RECT 7.905 1.755 8.335 2.125 ;
        RECT 6.535 1.495 7.725 1.665 ;
        RECT 5.105 0.885 5.410 0.925 ;
        RECT 7.470 0.885 7.775 0.925 ;
        RECT 8.025 0.885 8.195 1.755 ;
        RECT 8.550 1.645 8.720 2.295 ;
        RECT 8.990 1.635 9.320 2.465 ;
        RECT 8.890 1.475 9.320 1.635 ;
        RECT 8.540 1.465 9.320 1.475 ;
        RECT 9.495 1.465 9.825 2.635 ;
        RECT 10.000 1.635 10.330 2.465 ;
        RECT 10.600 2.295 11.765 2.465 ;
        RECT 10.600 1.645 10.770 2.295 ;
        RECT 10.985 1.755 11.415 2.125 ;
        RECT 10.000 1.475 10.430 1.635 ;
        RECT 10.000 1.465 10.780 1.475 ;
        RECT 8.540 1.305 9.060 1.465 ;
        RECT 10.260 1.305 10.780 1.465 ;
        RECT 8.540 1.205 8.955 1.305 ;
        RECT 2.345 0.585 2.925 0.755 ;
        RECT 1.030 0.255 2.175 0.425 ;
        RECT 2.675 0.330 2.925 0.585 ;
        RECT 3.095 0.085 3.345 0.660 ;
        RECT 3.515 0.585 4.095 0.755 ;
        RECT 3.515 0.330 3.765 0.585 ;
        RECT 4.265 0.425 4.435 0.770 ;
        RECT 4.605 0.595 4.935 0.885 ;
        RECT 5.105 0.715 6.295 0.885 ;
        RECT 5.105 0.425 5.410 0.715 ;
        RECT 4.265 0.255 5.410 0.425 ;
        RECT 5.580 0.085 5.795 0.545 ;
        RECT 5.965 0.255 6.295 0.715 ;
        RECT 6.585 0.715 7.775 0.885 ;
        RECT 6.585 0.255 6.915 0.715 ;
        RECT 7.085 0.085 7.300 0.545 ;
        RECT 7.470 0.425 7.775 0.715 ;
        RECT 7.945 0.595 8.275 0.885 ;
        RECT 8.445 0.425 8.615 0.770 ;
        RECT 8.785 0.755 8.955 1.205 ;
        RECT 10.365 1.205 10.780 1.305 ;
        RECT 10.365 0.755 10.535 1.205 ;
        RECT 11.125 0.885 11.295 1.755 ;
        RECT 11.595 1.665 11.765 2.295 ;
        RECT 11.985 2.105 12.285 2.635 ;
        RECT 12.455 2.210 12.785 2.465 ;
        RECT 11.985 1.835 12.315 2.105 ;
        RECT 12.485 1.665 12.785 2.210 ;
        RECT 11.595 1.495 12.785 1.665 ;
        RECT 11.545 0.885 11.850 0.925 ;
        RECT 8.785 0.585 9.365 0.755 ;
        RECT 7.470 0.255 8.615 0.425 ;
        RECT 9.115 0.330 9.365 0.585 ;
        RECT 9.535 0.085 9.785 0.660 ;
        RECT 9.955 0.585 10.535 0.755 ;
        RECT 9.955 0.330 10.205 0.585 ;
        RECT 10.705 0.425 10.875 0.770 ;
        RECT 11.045 0.595 11.375 0.885 ;
        RECT 11.545 0.715 12.735 0.885 ;
        RECT 11.545 0.425 11.850 0.715 ;
        RECT 10.705 0.255 11.850 0.425 ;
        RECT 12.020 0.085 12.235 0.545 ;
        RECT 12.405 0.255 12.735 0.715 ;
        RECT 0.000 -0.085 12.880 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 1.525 1.785 1.695 1.955 ;
        RECT 4.745 1.785 4.915 1.955 ;
        RECT 7.965 1.785 8.135 1.955 ;
        RECT 11.185 1.785 11.355 1.955 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__muxb4to1_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__muxb4to1_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__muxb4to1_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 23.975 1.055 25.365 1.325 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 13.275 1.055 14.665 1.325 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 11.095 1.055 12.485 1.325 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.395 1.055 1.785 1.325 ;
    END
  END D[0]
  PIN S[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.733200 ;
    PORT
      LAYER li1 ;
        RECT 19.405 0.995 20.000 1.325 ;
    END
  END S[3]
  PIN S[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.733200 ;
    PORT
      LAYER li1 ;
        RECT 18.640 0.995 19.235 1.325 ;
    END
  END S[2]
  PIN S[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.733200 ;
    PORT
      LAYER li1 ;
        RECT 6.525 0.995 7.120 1.325 ;
    END
  END S[1]
  PIN S[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.733200 ;
    PORT
      LAYER li1 ;
        RECT 5.760 0.995 6.355 1.325 ;
    END
  END S[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 25.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.980 2.345 1.015 ;
        RECT 10.535 0.980 15.225 1.015 ;
        RECT 23.415 0.980 25.755 1.015 ;
        RECT 0.005 0.785 4.545 0.980 ;
        RECT 8.335 0.785 17.425 0.980 ;
        RECT 21.215 0.785 25.755 0.980 ;
        RECT 0.005 0.200 25.755 0.785 ;
        RECT 0.005 0.105 2.345 0.200 ;
        RECT 4.910 0.105 7.970 0.200 ;
        RECT 10.535 0.105 15.225 0.200 ;
        RECT 17.790 0.105 20.850 0.200 ;
        RECT 23.415 0.105 25.755 0.200 ;
        RECT 0.145 -0.085 0.315 0.105 ;
        RECT 12.565 -0.085 13.195 0.105 ;
        RECT 25.445 -0.085 25.615 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 25.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 25.760 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.025600 ;
    PORT
      LAYER met1 ;
        RECT 2.985 1.940 3.275 1.985 ;
        RECT 3.925 1.940 4.215 1.985 ;
        RECT 8.665 1.940 8.955 1.985 ;
        RECT 9.605 1.940 9.895 1.985 ;
        RECT 15.865 1.940 16.155 1.985 ;
        RECT 16.805 1.940 17.095 1.985 ;
        RECT 21.545 1.940 21.835 1.985 ;
        RECT 22.485 1.940 22.775 1.985 ;
        RECT 2.985 1.800 22.775 1.940 ;
        RECT 2.985 1.755 3.275 1.800 ;
        RECT 3.925 1.755 4.215 1.800 ;
        RECT 8.665 1.755 8.955 1.800 ;
        RECT 9.605 1.755 9.895 1.800 ;
        RECT 15.865 1.755 16.155 1.800 ;
        RECT 16.805 1.755 17.095 1.800 ;
        RECT 21.545 1.755 21.835 1.800 ;
        RECT 22.485 1.755 22.775 1.800 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 25.760 2.805 ;
        RECT 0.125 1.495 0.395 2.635 ;
        RECT 0.565 1.665 0.895 2.465 ;
        RECT 1.065 1.835 1.335 2.635 ;
        RECT 1.505 1.665 1.835 2.465 ;
        RECT 2.005 1.835 2.275 2.635 ;
        RECT 2.495 2.295 4.705 2.465 ;
        RECT 2.495 1.665 2.795 2.295 ;
        RECT 0.565 1.495 2.795 1.665 ;
        RECT 2.965 1.365 3.295 2.125 ;
        RECT 3.465 1.535 3.735 2.295 ;
        RECT 3.905 1.365 4.235 2.125 ;
        RECT 4.405 1.565 4.705 2.295 ;
        RECT 4.950 1.605 5.225 2.635 ;
        RECT 5.420 1.605 5.750 2.465 ;
        RECT 5.920 1.605 6.220 2.635 ;
        RECT 6.660 1.605 6.960 2.635 ;
        RECT 7.130 1.605 7.460 2.465 ;
        RECT 7.655 1.605 7.930 2.635 ;
        RECT 8.175 2.295 10.385 2.465 ;
        RECT 5.420 1.395 5.590 1.605 ;
        RECT 2.965 1.065 4.235 1.365 ;
        RECT 4.405 1.065 5.590 1.395 ;
        RECT 2.965 0.885 3.195 1.065 ;
        RECT 0.145 0.085 0.395 0.885 ;
        RECT 0.565 0.715 2.695 0.885 ;
        RECT 0.565 0.255 0.895 0.715 ;
        RECT 1.065 0.085 1.335 0.545 ;
        RECT 1.505 0.255 1.835 0.715 ;
        RECT 2.005 0.085 2.255 0.545 ;
        RECT 2.425 0.425 2.695 0.715 ;
        RECT 2.865 0.595 3.195 0.885 ;
        RECT 3.365 0.425 3.535 0.770 ;
        RECT 3.705 0.595 4.035 1.065 ;
        RECT 5.420 0.825 5.590 1.065 ;
        RECT 7.290 1.395 7.460 1.605 ;
        RECT 8.175 1.565 8.475 2.295 ;
        RECT 7.290 1.065 8.475 1.395 ;
        RECT 8.645 1.365 8.975 2.125 ;
        RECT 9.145 1.535 9.415 2.295 ;
        RECT 9.585 1.365 9.915 2.125 ;
        RECT 10.085 1.665 10.385 2.295 ;
        RECT 10.605 1.835 10.875 2.635 ;
        RECT 11.045 1.665 11.375 2.465 ;
        RECT 11.545 1.835 11.815 2.635 ;
        RECT 11.985 1.665 12.315 2.465 ;
        RECT 10.085 1.495 12.315 1.665 ;
        RECT 12.485 1.495 12.755 2.635 ;
        RECT 13.005 1.495 13.275 2.635 ;
        RECT 13.445 1.665 13.775 2.465 ;
        RECT 13.945 1.835 14.215 2.635 ;
        RECT 14.385 1.665 14.715 2.465 ;
        RECT 14.885 1.835 15.155 2.635 ;
        RECT 15.375 2.295 17.585 2.465 ;
        RECT 15.375 1.665 15.675 2.295 ;
        RECT 13.445 1.495 15.675 1.665 ;
        RECT 8.645 1.065 9.915 1.365 ;
        RECT 7.290 0.825 7.460 1.065 ;
        RECT 4.205 0.425 4.455 0.770 ;
        RECT 2.425 0.255 4.455 0.425 ;
        RECT 4.960 0.085 5.250 0.610 ;
        RECT 5.420 0.280 5.670 0.825 ;
        RECT 5.880 0.085 6.170 0.610 ;
        RECT 6.710 0.085 7.000 0.610 ;
        RECT 7.210 0.280 7.460 0.825 ;
        RECT 7.630 0.085 7.920 0.610 ;
        RECT 8.425 0.425 8.675 0.770 ;
        RECT 8.845 0.595 9.175 1.065 ;
        RECT 9.685 0.885 9.915 1.065 ;
        RECT 15.845 1.365 16.175 2.125 ;
        RECT 16.345 1.535 16.615 2.295 ;
        RECT 16.785 1.365 17.115 2.125 ;
        RECT 17.285 1.565 17.585 2.295 ;
        RECT 17.830 1.605 18.105 2.635 ;
        RECT 18.300 1.605 18.630 2.465 ;
        RECT 18.800 1.605 19.100 2.635 ;
        RECT 19.540 1.605 19.840 2.635 ;
        RECT 20.010 1.605 20.340 2.465 ;
        RECT 20.535 1.605 20.810 2.635 ;
        RECT 21.055 2.295 23.265 2.465 ;
        RECT 18.300 1.395 18.470 1.605 ;
        RECT 15.845 1.065 17.115 1.365 ;
        RECT 17.285 1.065 18.470 1.395 ;
        RECT 15.845 0.885 16.075 1.065 ;
        RECT 9.345 0.425 9.515 0.770 ;
        RECT 9.685 0.595 10.015 0.885 ;
        RECT 10.185 0.715 12.315 0.885 ;
        RECT 10.185 0.425 10.455 0.715 ;
        RECT 8.425 0.255 10.455 0.425 ;
        RECT 10.625 0.085 10.875 0.545 ;
        RECT 11.045 0.255 11.375 0.715 ;
        RECT 11.545 0.085 11.815 0.545 ;
        RECT 11.985 0.255 12.315 0.715 ;
        RECT 12.485 0.085 12.735 0.885 ;
        RECT 13.025 0.085 13.275 0.885 ;
        RECT 13.445 0.715 15.575 0.885 ;
        RECT 13.445 0.255 13.775 0.715 ;
        RECT 13.945 0.085 14.215 0.545 ;
        RECT 14.385 0.255 14.715 0.715 ;
        RECT 14.885 0.085 15.135 0.545 ;
        RECT 15.305 0.425 15.575 0.715 ;
        RECT 15.745 0.595 16.075 0.885 ;
        RECT 16.245 0.425 16.415 0.770 ;
        RECT 16.585 0.595 16.915 1.065 ;
        RECT 18.300 0.825 18.470 1.065 ;
        RECT 20.170 1.395 20.340 1.605 ;
        RECT 21.055 1.565 21.355 2.295 ;
        RECT 20.170 1.065 21.355 1.395 ;
        RECT 21.525 1.365 21.855 2.125 ;
        RECT 22.025 1.535 22.295 2.295 ;
        RECT 22.465 1.365 22.795 2.125 ;
        RECT 22.965 1.665 23.265 2.295 ;
        RECT 23.485 1.835 23.755 2.635 ;
        RECT 23.925 1.665 24.255 2.465 ;
        RECT 24.425 1.835 24.695 2.635 ;
        RECT 24.865 1.665 25.195 2.465 ;
        RECT 22.965 1.495 25.195 1.665 ;
        RECT 25.365 1.495 25.635 2.635 ;
        RECT 21.525 1.065 22.795 1.365 ;
        RECT 20.170 0.825 20.340 1.065 ;
        RECT 17.085 0.425 17.335 0.770 ;
        RECT 15.305 0.255 17.335 0.425 ;
        RECT 17.840 0.085 18.130 0.610 ;
        RECT 18.300 0.280 18.550 0.825 ;
        RECT 18.760 0.085 19.050 0.610 ;
        RECT 19.590 0.085 19.880 0.610 ;
        RECT 20.090 0.280 20.340 0.825 ;
        RECT 20.510 0.085 20.800 0.610 ;
        RECT 21.305 0.425 21.555 0.770 ;
        RECT 21.725 0.595 22.055 1.065 ;
        RECT 22.565 0.885 22.795 1.065 ;
        RECT 22.225 0.425 22.395 0.770 ;
        RECT 22.565 0.595 22.895 0.885 ;
        RECT 23.065 0.715 25.195 0.885 ;
        RECT 23.065 0.425 23.335 0.715 ;
        RECT 21.305 0.255 23.335 0.425 ;
        RECT 23.505 0.085 23.755 0.545 ;
        RECT 23.925 0.255 24.255 0.715 ;
        RECT 24.425 0.085 24.695 0.545 ;
        RECT 24.865 0.255 25.195 0.715 ;
        RECT 25.365 0.085 25.615 0.885 ;
        RECT 0.000 -0.085 25.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 14.405 2.635 14.575 2.805 ;
        RECT 14.865 2.635 15.035 2.805 ;
        RECT 15.325 2.635 15.495 2.805 ;
        RECT 15.785 2.635 15.955 2.805 ;
        RECT 16.245 2.635 16.415 2.805 ;
        RECT 16.705 2.635 16.875 2.805 ;
        RECT 17.165 2.635 17.335 2.805 ;
        RECT 17.625 2.635 17.795 2.805 ;
        RECT 18.085 2.635 18.255 2.805 ;
        RECT 18.545 2.635 18.715 2.805 ;
        RECT 19.005 2.635 19.175 2.805 ;
        RECT 19.465 2.635 19.635 2.805 ;
        RECT 19.925 2.635 20.095 2.805 ;
        RECT 20.385 2.635 20.555 2.805 ;
        RECT 20.845 2.635 21.015 2.805 ;
        RECT 21.305 2.635 21.475 2.805 ;
        RECT 21.765 2.635 21.935 2.805 ;
        RECT 22.225 2.635 22.395 2.805 ;
        RECT 22.685 2.635 22.855 2.805 ;
        RECT 23.145 2.635 23.315 2.805 ;
        RECT 23.605 2.635 23.775 2.805 ;
        RECT 24.065 2.635 24.235 2.805 ;
        RECT 24.525 2.635 24.695 2.805 ;
        RECT 24.985 2.635 25.155 2.805 ;
        RECT 25.445 2.635 25.615 2.805 ;
        RECT 3.045 1.785 3.215 1.955 ;
        RECT 3.985 1.785 4.155 1.955 ;
        RECT 8.725 1.785 8.895 1.955 ;
        RECT 9.665 1.785 9.835 1.955 ;
        RECT 15.925 1.785 16.095 1.955 ;
        RECT 16.865 1.785 17.035 1.955 ;
        RECT 21.605 1.785 21.775 1.955 ;
        RECT 22.545 1.785 22.715 1.955 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
        RECT 14.405 -0.085 14.575 0.085 ;
        RECT 14.865 -0.085 15.035 0.085 ;
        RECT 15.325 -0.085 15.495 0.085 ;
        RECT 15.785 -0.085 15.955 0.085 ;
        RECT 16.245 -0.085 16.415 0.085 ;
        RECT 16.705 -0.085 16.875 0.085 ;
        RECT 17.165 -0.085 17.335 0.085 ;
        RECT 17.625 -0.085 17.795 0.085 ;
        RECT 18.085 -0.085 18.255 0.085 ;
        RECT 18.545 -0.085 18.715 0.085 ;
        RECT 19.005 -0.085 19.175 0.085 ;
        RECT 19.465 -0.085 19.635 0.085 ;
        RECT 19.925 -0.085 20.095 0.085 ;
        RECT 20.385 -0.085 20.555 0.085 ;
        RECT 20.845 -0.085 21.015 0.085 ;
        RECT 21.305 -0.085 21.475 0.085 ;
        RECT 21.765 -0.085 21.935 0.085 ;
        RECT 22.225 -0.085 22.395 0.085 ;
        RECT 22.685 -0.085 22.855 0.085 ;
        RECT 23.145 -0.085 23.315 0.085 ;
        RECT 23.605 -0.085 23.775 0.085 ;
        RECT 24.065 -0.085 24.235 0.085 ;
        RECT 24.525 -0.085 24.695 0.085 ;
        RECT 24.985 -0.085 25.155 0.085 ;
        RECT 25.445 -0.085 25.615 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__muxb4to1_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__muxb8to1_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__muxb8to1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.020 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 16.290 1.055 16.685 1.325 ;
        RECT 16.290 0.625 16.460 1.055 ;
        RECT 16.185 0.395 16.460 0.625 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 12.755 1.055 13.150 1.325 ;
        RECT 12.980 0.625 13.150 1.055 ;
        RECT 12.980 0.395 13.255 0.625 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 12.150 1.055 12.545 1.325 ;
        RECT 12.150 0.625 12.320 1.055 ;
        RECT 12.045 0.395 12.320 0.625 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 8.615 1.055 9.010 1.325 ;
        RECT 8.840 0.625 9.010 1.055 ;
        RECT 8.840 0.395 9.115 0.625 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 8.010 1.055 8.405 1.325 ;
        RECT 8.010 0.625 8.180 1.055 ;
        RECT 7.905 0.395 8.180 0.625 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 4.475 1.055 4.870 1.325 ;
        RECT 4.700 0.625 4.870 1.055 ;
        RECT 4.700 0.395 4.975 0.625 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 3.870 1.055 4.265 1.325 ;
        RECT 3.870 0.625 4.040 1.055 ;
        RECT 3.765 0.395 4.040 0.625 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.335 1.055 0.730 1.325 ;
        RECT 0.560 0.625 0.730 1.055 ;
        RECT 0.560 0.395 0.835 0.625 ;
    END
  END D[0]
  PIN S[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 14.815 0.945 15.215 1.295 ;
    END
  END S[7]
  PIN S[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 14.225 0.945 14.625 1.295 ;
    END
  END S[6]
  PIN S[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 10.675 0.945 11.075 1.295 ;
    END
  END S[5]
  PIN S[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 10.085 0.945 10.485 1.295 ;
    END
  END S[4]
  PIN S[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 6.535 0.945 6.935 1.295 ;
    END
  END S[3]
  PIN S[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 5.945 0.945 6.345 1.295 ;
    END
  END S[2]
  PIN S[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 2.395 0.945 2.795 1.295 ;
    END
  END S[1]
  PIN S[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 1.805 0.945 2.205 1.295 ;
    END
  END S[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 17.020 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.885 0.925 1.015 ;
        RECT 3.675 0.885 5.065 1.015 ;
        RECT 7.815 0.885 9.205 1.015 ;
        RECT 11.955 0.885 13.345 1.015 ;
        RECT 16.095 0.885 17.015 1.015 ;
        RECT 0.005 0.105 17.015 0.885 ;
        RECT 0.145 -0.085 0.315 0.105 ;
        RECT 4.285 -0.085 4.455 0.105 ;
        RECT 8.425 -0.085 8.595 0.105 ;
        RECT 12.565 -0.085 12.735 0.105 ;
        RECT 16.705 -0.085 16.875 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 17.210 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 17.020 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.852800 ;
    PORT
      LAYER met1 ;
        RECT 1.005 1.940 1.295 1.985 ;
        RECT 3.305 1.940 3.595 1.985 ;
        RECT 5.145 1.940 5.435 1.985 ;
        RECT 7.445 1.940 7.735 1.985 ;
        RECT 9.285 1.940 9.575 1.985 ;
        RECT 11.585 1.940 11.875 1.985 ;
        RECT 13.425 1.940 13.715 1.985 ;
        RECT 15.725 1.940 16.015 1.985 ;
        RECT 1.005 1.800 16.015 1.940 ;
        RECT 1.005 1.755 1.295 1.800 ;
        RECT 3.305 1.755 3.595 1.800 ;
        RECT 5.145 1.755 5.435 1.800 ;
        RECT 7.445 1.755 7.735 1.800 ;
        RECT 9.285 1.755 9.575 1.800 ;
        RECT 11.585 1.755 11.875 1.800 ;
        RECT 13.425 1.755 13.715 1.800 ;
        RECT 15.725 1.755 16.015 1.800 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 17.020 2.805 ;
        RECT 0.095 1.495 0.425 2.635 ;
        RECT 1.090 1.985 1.420 2.465 ;
        RECT 0.900 1.805 1.420 1.985 ;
        RECT 0.900 1.755 1.295 1.805 ;
        RECT 0.900 1.005 1.070 1.755 ;
        RECT 1.610 1.635 1.940 2.465 ;
        RECT 1.460 1.505 1.940 1.635 ;
        RECT 1.240 1.465 1.940 1.505 ;
        RECT 2.135 1.465 2.465 2.635 ;
        RECT 2.660 1.635 2.990 2.465 ;
        RECT 3.180 1.985 3.510 2.465 ;
        RECT 3.180 1.805 3.700 1.985 ;
        RECT 3.305 1.755 3.700 1.805 ;
        RECT 2.660 1.505 3.140 1.635 ;
        RECT 2.660 1.465 3.360 1.505 ;
        RECT 1.240 1.175 1.630 1.465 ;
        RECT 0.130 0.085 0.390 0.885 ;
        RECT 0.900 0.835 1.290 1.005 ;
        RECT 1.045 0.330 1.290 0.835 ;
        RECT 1.460 0.755 1.630 1.175 ;
        RECT 2.970 1.175 3.360 1.465 ;
        RECT 2.970 0.755 3.140 1.175 ;
        RECT 3.530 1.005 3.700 1.755 ;
        RECT 4.175 1.495 4.565 2.635 ;
        RECT 5.230 1.985 5.560 2.465 ;
        RECT 5.040 1.805 5.560 1.985 ;
        RECT 5.040 1.755 5.435 1.805 ;
        RECT 1.460 0.585 1.900 0.755 ;
        RECT 1.650 0.330 1.900 0.585 ;
        RECT 2.135 0.085 2.465 0.660 ;
        RECT 2.700 0.585 3.140 0.755 ;
        RECT 3.310 0.835 3.700 1.005 ;
        RECT 5.040 1.005 5.210 1.755 ;
        RECT 5.750 1.635 6.080 2.465 ;
        RECT 5.600 1.505 6.080 1.635 ;
        RECT 5.380 1.465 6.080 1.505 ;
        RECT 6.275 1.465 6.605 2.635 ;
        RECT 6.800 1.635 7.130 2.465 ;
        RECT 7.320 1.985 7.650 2.465 ;
        RECT 7.320 1.805 7.840 1.985 ;
        RECT 7.445 1.755 7.840 1.805 ;
        RECT 6.800 1.505 7.280 1.635 ;
        RECT 6.800 1.465 7.500 1.505 ;
        RECT 5.380 1.175 5.770 1.465 ;
        RECT 2.700 0.330 2.950 0.585 ;
        RECT 3.310 0.330 3.555 0.835 ;
        RECT 4.210 0.085 4.530 0.885 ;
        RECT 5.040 0.835 5.430 1.005 ;
        RECT 5.185 0.330 5.430 0.835 ;
        RECT 5.600 0.755 5.770 1.175 ;
        RECT 7.110 1.175 7.500 1.465 ;
        RECT 7.110 0.755 7.280 1.175 ;
        RECT 7.670 1.005 7.840 1.755 ;
        RECT 8.315 1.495 8.705 2.635 ;
        RECT 9.370 1.985 9.700 2.465 ;
        RECT 9.180 1.805 9.700 1.985 ;
        RECT 9.180 1.755 9.575 1.805 ;
        RECT 5.600 0.585 6.040 0.755 ;
        RECT 5.790 0.330 6.040 0.585 ;
        RECT 6.275 0.085 6.605 0.660 ;
        RECT 6.840 0.585 7.280 0.755 ;
        RECT 7.450 0.835 7.840 1.005 ;
        RECT 9.180 1.005 9.350 1.755 ;
        RECT 9.890 1.635 10.220 2.465 ;
        RECT 9.740 1.505 10.220 1.635 ;
        RECT 9.520 1.465 10.220 1.505 ;
        RECT 10.415 1.465 10.745 2.635 ;
        RECT 10.940 1.635 11.270 2.465 ;
        RECT 11.460 1.985 11.790 2.465 ;
        RECT 11.460 1.805 11.980 1.985 ;
        RECT 11.585 1.755 11.980 1.805 ;
        RECT 10.940 1.505 11.420 1.635 ;
        RECT 10.940 1.465 11.640 1.505 ;
        RECT 9.520 1.175 9.910 1.465 ;
        RECT 6.840 0.330 7.090 0.585 ;
        RECT 7.450 0.330 7.695 0.835 ;
        RECT 8.350 0.085 8.670 0.885 ;
        RECT 9.180 0.835 9.570 1.005 ;
        RECT 9.325 0.330 9.570 0.835 ;
        RECT 9.740 0.755 9.910 1.175 ;
        RECT 11.250 1.175 11.640 1.465 ;
        RECT 11.250 0.755 11.420 1.175 ;
        RECT 11.810 1.005 11.980 1.755 ;
        RECT 12.455 1.495 12.845 2.635 ;
        RECT 13.510 1.985 13.840 2.465 ;
        RECT 13.320 1.805 13.840 1.985 ;
        RECT 13.320 1.755 13.715 1.805 ;
        RECT 9.740 0.585 10.180 0.755 ;
        RECT 9.930 0.330 10.180 0.585 ;
        RECT 10.415 0.085 10.745 0.660 ;
        RECT 10.980 0.585 11.420 0.755 ;
        RECT 11.590 0.835 11.980 1.005 ;
        RECT 13.320 1.005 13.490 1.755 ;
        RECT 14.030 1.635 14.360 2.465 ;
        RECT 13.880 1.505 14.360 1.635 ;
        RECT 13.660 1.465 14.360 1.505 ;
        RECT 14.555 1.465 14.885 2.635 ;
        RECT 15.080 1.635 15.410 2.465 ;
        RECT 15.600 1.985 15.930 2.465 ;
        RECT 15.600 1.805 16.120 1.985 ;
        RECT 15.725 1.755 16.120 1.805 ;
        RECT 15.080 1.505 15.560 1.635 ;
        RECT 15.080 1.465 15.780 1.505 ;
        RECT 13.660 1.175 14.050 1.465 ;
        RECT 10.980 0.330 11.230 0.585 ;
        RECT 11.590 0.330 11.835 0.835 ;
        RECT 12.490 0.085 12.810 0.885 ;
        RECT 13.320 0.835 13.710 1.005 ;
        RECT 13.465 0.330 13.710 0.835 ;
        RECT 13.880 0.755 14.050 1.175 ;
        RECT 15.390 1.175 15.780 1.465 ;
        RECT 15.390 0.755 15.560 1.175 ;
        RECT 15.950 1.005 16.120 1.755 ;
        RECT 16.595 1.495 16.925 2.635 ;
        RECT 13.880 0.585 14.320 0.755 ;
        RECT 14.070 0.330 14.320 0.585 ;
        RECT 14.555 0.085 14.885 0.660 ;
        RECT 15.120 0.585 15.560 0.755 ;
        RECT 15.730 0.835 16.120 1.005 ;
        RECT 15.120 0.330 15.370 0.585 ;
        RECT 15.730 0.330 15.975 0.835 ;
        RECT 16.630 0.085 16.890 0.885 ;
        RECT 0.000 -0.085 17.020 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 14.405 2.635 14.575 2.805 ;
        RECT 14.865 2.635 15.035 2.805 ;
        RECT 15.325 2.635 15.495 2.805 ;
        RECT 15.785 2.635 15.955 2.805 ;
        RECT 16.245 2.635 16.415 2.805 ;
        RECT 16.705 2.635 16.875 2.805 ;
        RECT 1.065 1.785 1.235 1.955 ;
        RECT 3.365 1.785 3.535 1.955 ;
        RECT 5.205 1.785 5.375 1.955 ;
        RECT 7.505 1.785 7.675 1.955 ;
        RECT 9.345 1.785 9.515 1.955 ;
        RECT 11.645 1.785 11.815 1.955 ;
        RECT 13.485 1.785 13.655 1.955 ;
        RECT 15.785 1.785 15.955 1.955 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
        RECT 14.405 -0.085 14.575 0.085 ;
        RECT 14.865 -0.085 15.035 0.085 ;
        RECT 15.325 -0.085 15.495 0.085 ;
        RECT 15.785 -0.085 15.955 0.085 ;
        RECT 16.245 -0.085 16.415 0.085 ;
        RECT 16.705 -0.085 16.875 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__muxb8to1_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__muxb8to1_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__muxb8to1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 24.845 1.055 25.665 1.325 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 19.415 1.055 20.235 1.325 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 18.405 1.055 19.225 1.325 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 12.975 1.055 13.795 1.325 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 11.965 1.055 12.785 1.325 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 6.535 1.055 7.355 1.325 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 5.525 1.055 6.345 1.325 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.055 0.915 1.325 ;
    END
  END D[0]
  PIN S[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 22.635 1.025 22.970 1.295 ;
    END
  END S[7]
  PIN S[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 22.110 1.025 22.445 1.295 ;
    END
  END S[6]
  PIN S[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 16.195 1.025 16.530 1.295 ;
    END
  END S[5]
  PIN S[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 15.670 1.025 16.005 1.295 ;
    END
  END S[4]
  PIN S[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 9.755 1.025 10.090 1.295 ;
    END
  END S[3]
  PIN S[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 9.230 1.025 9.565 1.295 ;
    END
  END S[2]
  PIN S[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 3.315 1.025 3.650 1.295 ;
    END
  END S[1]
  PIN S[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 2.790 1.025 3.125 1.295 ;
    END
  END S[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 25.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.995 1.440 1.015 ;
        RECT 5.000 0.995 7.880 1.015 ;
        RECT 11.440 0.995 14.320 1.015 ;
        RECT 17.880 0.995 20.760 1.015 ;
        RECT 24.320 0.995 25.755 1.015 ;
        RECT 0.005 0.885 2.345 0.995 ;
        RECT 4.095 0.885 8.785 0.995 ;
        RECT 10.535 0.885 15.225 0.995 ;
        RECT 16.975 0.885 21.665 0.995 ;
        RECT 23.415 0.885 25.755 0.995 ;
        RECT 0.005 0.215 25.755 0.885 ;
        RECT 0.005 0.105 1.440 0.215 ;
        RECT 2.545 0.105 3.895 0.215 ;
        RECT 5.000 0.105 7.880 0.215 ;
        RECT 8.985 0.105 10.335 0.215 ;
        RECT 11.440 0.105 14.320 0.215 ;
        RECT 15.425 0.105 16.775 0.215 ;
        RECT 17.880 0.105 20.760 0.215 ;
        RECT 21.865 0.105 23.215 0.215 ;
        RECT 24.320 0.105 25.755 0.215 ;
        RECT 0.145 -0.085 0.315 0.105 ;
        RECT 6.125 -0.085 6.755 0.105 ;
        RECT 12.565 -0.085 13.195 0.105 ;
        RECT 19.005 -0.085 19.635 0.105 ;
        RECT 25.445 -0.085 25.615 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 25.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 25.760 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.025600 ;
    PORT
      LAYER met1 ;
        RECT 1.465 1.940 1.755 1.985 ;
        RECT 4.685 1.940 4.975 1.985 ;
        RECT 7.905 1.940 8.195 1.985 ;
        RECT 11.125 1.940 11.415 1.985 ;
        RECT 14.345 1.940 14.635 1.985 ;
        RECT 17.565 1.940 17.855 1.985 ;
        RECT 20.785 1.940 21.075 1.985 ;
        RECT 24.005 1.940 24.295 1.985 ;
        RECT 1.465 1.800 24.295 1.940 ;
        RECT 1.465 1.755 1.755 1.800 ;
        RECT 4.685 1.755 4.975 1.800 ;
        RECT 7.905 1.755 8.195 1.800 ;
        RECT 11.125 1.755 11.415 1.800 ;
        RECT 14.345 1.755 14.635 1.800 ;
        RECT 17.565 1.755 17.855 1.800 ;
        RECT 20.785 1.755 21.075 1.800 ;
        RECT 24.005 1.755 24.295 1.800 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 25.760 2.805 ;
        RECT 0.095 2.210 0.425 2.465 ;
        RECT 0.095 1.665 0.395 2.210 ;
        RECT 0.595 2.105 0.895 2.635 ;
        RECT 0.565 1.835 0.895 2.105 ;
        RECT 1.115 2.295 2.280 2.465 ;
        RECT 1.115 1.665 1.285 2.295 ;
        RECT 1.465 1.755 1.895 2.125 ;
        RECT 0.095 1.495 1.285 1.665 ;
        RECT 1.030 0.885 1.335 0.925 ;
        RECT 1.585 0.885 1.755 1.755 ;
        RECT 2.110 1.645 2.280 2.295 ;
        RECT 2.550 1.635 2.880 2.465 ;
        RECT 2.450 1.475 2.880 1.635 ;
        RECT 2.100 1.465 2.880 1.475 ;
        RECT 3.055 1.465 3.385 2.635 ;
        RECT 3.560 1.635 3.890 2.465 ;
        RECT 4.160 2.295 5.325 2.465 ;
        RECT 4.160 1.645 4.330 2.295 ;
        RECT 4.545 1.755 4.975 2.125 ;
        RECT 3.560 1.475 3.990 1.635 ;
        RECT 3.560 1.465 4.340 1.475 ;
        RECT 2.100 1.305 2.620 1.465 ;
        RECT 3.820 1.305 4.340 1.465 ;
        RECT 2.100 1.205 2.515 1.305 ;
        RECT 0.145 0.715 1.335 0.885 ;
        RECT 0.145 0.255 0.475 0.715 ;
        RECT 0.645 0.085 0.860 0.545 ;
        RECT 1.030 0.425 1.335 0.715 ;
        RECT 1.505 0.595 1.835 0.885 ;
        RECT 2.005 0.425 2.175 0.770 ;
        RECT 2.345 0.755 2.515 1.205 ;
        RECT 3.925 1.205 4.340 1.305 ;
        RECT 3.925 0.755 4.095 1.205 ;
        RECT 4.685 0.885 4.855 1.755 ;
        RECT 5.155 1.665 5.325 2.295 ;
        RECT 5.545 2.105 5.845 2.635 ;
        RECT 6.015 2.210 6.345 2.465 ;
        RECT 5.545 1.835 5.875 2.105 ;
        RECT 6.045 1.665 6.345 2.210 ;
        RECT 5.155 1.495 6.345 1.665 ;
        RECT 6.535 2.210 6.865 2.465 ;
        RECT 6.535 1.665 6.835 2.210 ;
        RECT 7.035 2.105 7.335 2.635 ;
        RECT 7.005 1.835 7.335 2.105 ;
        RECT 7.555 2.295 8.720 2.465 ;
        RECT 7.555 1.665 7.725 2.295 ;
        RECT 7.905 1.755 8.335 2.125 ;
        RECT 6.535 1.495 7.725 1.665 ;
        RECT 5.105 0.885 5.410 0.925 ;
        RECT 7.470 0.885 7.775 0.925 ;
        RECT 8.025 0.885 8.195 1.755 ;
        RECT 8.550 1.645 8.720 2.295 ;
        RECT 8.990 1.635 9.320 2.465 ;
        RECT 8.890 1.475 9.320 1.635 ;
        RECT 8.540 1.465 9.320 1.475 ;
        RECT 9.495 1.465 9.825 2.635 ;
        RECT 10.000 1.635 10.330 2.465 ;
        RECT 10.600 2.295 11.765 2.465 ;
        RECT 10.600 1.645 10.770 2.295 ;
        RECT 10.985 1.755 11.415 2.125 ;
        RECT 10.000 1.475 10.430 1.635 ;
        RECT 10.000 1.465 10.780 1.475 ;
        RECT 8.540 1.305 9.060 1.465 ;
        RECT 10.260 1.305 10.780 1.465 ;
        RECT 8.540 1.205 8.955 1.305 ;
        RECT 2.345 0.585 2.925 0.755 ;
        RECT 1.030 0.255 2.175 0.425 ;
        RECT 2.675 0.330 2.925 0.585 ;
        RECT 3.095 0.085 3.345 0.660 ;
        RECT 3.515 0.585 4.095 0.755 ;
        RECT 3.515 0.330 3.765 0.585 ;
        RECT 4.265 0.425 4.435 0.770 ;
        RECT 4.605 0.595 4.935 0.885 ;
        RECT 5.105 0.715 6.295 0.885 ;
        RECT 5.105 0.425 5.410 0.715 ;
        RECT 4.265 0.255 5.410 0.425 ;
        RECT 5.580 0.085 5.795 0.545 ;
        RECT 5.965 0.255 6.295 0.715 ;
        RECT 6.585 0.715 7.775 0.885 ;
        RECT 6.585 0.255 6.915 0.715 ;
        RECT 7.085 0.085 7.300 0.545 ;
        RECT 7.470 0.425 7.775 0.715 ;
        RECT 7.945 0.595 8.275 0.885 ;
        RECT 8.445 0.425 8.615 0.770 ;
        RECT 8.785 0.755 8.955 1.205 ;
        RECT 10.365 1.205 10.780 1.305 ;
        RECT 10.365 0.755 10.535 1.205 ;
        RECT 11.125 0.885 11.295 1.755 ;
        RECT 11.595 1.665 11.765 2.295 ;
        RECT 11.985 2.105 12.285 2.635 ;
        RECT 12.455 2.210 12.785 2.465 ;
        RECT 11.985 1.835 12.315 2.105 ;
        RECT 12.485 1.665 12.785 2.210 ;
        RECT 11.595 1.495 12.785 1.665 ;
        RECT 12.975 2.210 13.305 2.465 ;
        RECT 12.975 1.665 13.275 2.210 ;
        RECT 13.475 2.105 13.775 2.635 ;
        RECT 13.445 1.835 13.775 2.105 ;
        RECT 13.995 2.295 15.160 2.465 ;
        RECT 13.995 1.665 14.165 2.295 ;
        RECT 14.345 1.755 14.775 2.125 ;
        RECT 12.975 1.495 14.165 1.665 ;
        RECT 11.545 0.885 11.850 0.925 ;
        RECT 13.910 0.885 14.215 0.925 ;
        RECT 14.465 0.885 14.635 1.755 ;
        RECT 14.990 1.645 15.160 2.295 ;
        RECT 15.430 1.635 15.760 2.465 ;
        RECT 15.330 1.475 15.760 1.635 ;
        RECT 14.980 1.465 15.760 1.475 ;
        RECT 15.935 1.465 16.265 2.635 ;
        RECT 16.440 1.635 16.770 2.465 ;
        RECT 17.040 2.295 18.205 2.465 ;
        RECT 17.040 1.645 17.210 2.295 ;
        RECT 17.425 1.755 17.855 2.125 ;
        RECT 16.440 1.475 16.870 1.635 ;
        RECT 16.440 1.465 17.220 1.475 ;
        RECT 14.980 1.305 15.500 1.465 ;
        RECT 16.700 1.305 17.220 1.465 ;
        RECT 14.980 1.205 15.395 1.305 ;
        RECT 8.785 0.585 9.365 0.755 ;
        RECT 7.470 0.255 8.615 0.425 ;
        RECT 9.115 0.330 9.365 0.585 ;
        RECT 9.535 0.085 9.785 0.660 ;
        RECT 9.955 0.585 10.535 0.755 ;
        RECT 9.955 0.330 10.205 0.585 ;
        RECT 10.705 0.425 10.875 0.770 ;
        RECT 11.045 0.595 11.375 0.885 ;
        RECT 11.545 0.715 12.735 0.885 ;
        RECT 11.545 0.425 11.850 0.715 ;
        RECT 10.705 0.255 11.850 0.425 ;
        RECT 12.020 0.085 12.235 0.545 ;
        RECT 12.405 0.255 12.735 0.715 ;
        RECT 13.025 0.715 14.215 0.885 ;
        RECT 13.025 0.255 13.355 0.715 ;
        RECT 13.525 0.085 13.740 0.545 ;
        RECT 13.910 0.425 14.215 0.715 ;
        RECT 14.385 0.595 14.715 0.885 ;
        RECT 14.885 0.425 15.055 0.770 ;
        RECT 15.225 0.755 15.395 1.205 ;
        RECT 16.805 1.205 17.220 1.305 ;
        RECT 16.805 0.755 16.975 1.205 ;
        RECT 17.565 0.885 17.735 1.755 ;
        RECT 18.035 1.665 18.205 2.295 ;
        RECT 18.425 2.105 18.725 2.635 ;
        RECT 18.895 2.210 19.225 2.465 ;
        RECT 18.425 1.835 18.755 2.105 ;
        RECT 18.925 1.665 19.225 2.210 ;
        RECT 18.035 1.495 19.225 1.665 ;
        RECT 19.415 2.210 19.745 2.465 ;
        RECT 19.415 1.665 19.715 2.210 ;
        RECT 19.915 2.105 20.215 2.635 ;
        RECT 19.885 1.835 20.215 2.105 ;
        RECT 20.435 2.295 21.600 2.465 ;
        RECT 20.435 1.665 20.605 2.295 ;
        RECT 20.785 1.755 21.215 2.125 ;
        RECT 19.415 1.495 20.605 1.665 ;
        RECT 17.985 0.885 18.290 0.925 ;
        RECT 20.350 0.885 20.655 0.925 ;
        RECT 20.905 0.885 21.075 1.755 ;
        RECT 21.430 1.645 21.600 2.295 ;
        RECT 21.870 1.635 22.200 2.465 ;
        RECT 21.770 1.475 22.200 1.635 ;
        RECT 21.420 1.465 22.200 1.475 ;
        RECT 22.375 1.465 22.705 2.635 ;
        RECT 22.880 1.635 23.210 2.465 ;
        RECT 23.480 2.295 24.645 2.465 ;
        RECT 23.480 1.645 23.650 2.295 ;
        RECT 23.865 1.755 24.295 2.125 ;
        RECT 22.880 1.475 23.310 1.635 ;
        RECT 22.880 1.465 23.660 1.475 ;
        RECT 21.420 1.305 21.940 1.465 ;
        RECT 23.140 1.305 23.660 1.465 ;
        RECT 21.420 1.205 21.835 1.305 ;
        RECT 15.225 0.585 15.805 0.755 ;
        RECT 13.910 0.255 15.055 0.425 ;
        RECT 15.555 0.330 15.805 0.585 ;
        RECT 15.975 0.085 16.225 0.660 ;
        RECT 16.395 0.585 16.975 0.755 ;
        RECT 16.395 0.330 16.645 0.585 ;
        RECT 17.145 0.425 17.315 0.770 ;
        RECT 17.485 0.595 17.815 0.885 ;
        RECT 17.985 0.715 19.175 0.885 ;
        RECT 17.985 0.425 18.290 0.715 ;
        RECT 17.145 0.255 18.290 0.425 ;
        RECT 18.460 0.085 18.675 0.545 ;
        RECT 18.845 0.255 19.175 0.715 ;
        RECT 19.465 0.715 20.655 0.885 ;
        RECT 19.465 0.255 19.795 0.715 ;
        RECT 19.965 0.085 20.180 0.545 ;
        RECT 20.350 0.425 20.655 0.715 ;
        RECT 20.825 0.595 21.155 0.885 ;
        RECT 21.325 0.425 21.495 0.770 ;
        RECT 21.665 0.755 21.835 1.205 ;
        RECT 23.245 1.205 23.660 1.305 ;
        RECT 23.245 0.755 23.415 1.205 ;
        RECT 24.005 0.885 24.175 1.755 ;
        RECT 24.475 1.665 24.645 2.295 ;
        RECT 24.865 2.105 25.165 2.635 ;
        RECT 25.335 2.210 25.665 2.465 ;
        RECT 24.865 1.835 25.195 2.105 ;
        RECT 25.365 1.665 25.665 2.210 ;
        RECT 24.475 1.495 25.665 1.665 ;
        RECT 24.425 0.885 24.730 0.925 ;
        RECT 21.665 0.585 22.245 0.755 ;
        RECT 20.350 0.255 21.495 0.425 ;
        RECT 21.995 0.330 22.245 0.585 ;
        RECT 22.415 0.085 22.665 0.660 ;
        RECT 22.835 0.585 23.415 0.755 ;
        RECT 22.835 0.330 23.085 0.585 ;
        RECT 23.585 0.425 23.755 0.770 ;
        RECT 23.925 0.595 24.255 0.885 ;
        RECT 24.425 0.715 25.615 0.885 ;
        RECT 24.425 0.425 24.730 0.715 ;
        RECT 23.585 0.255 24.730 0.425 ;
        RECT 24.900 0.085 25.115 0.545 ;
        RECT 25.285 0.255 25.615 0.715 ;
        RECT 0.000 -0.085 25.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 14.405 2.635 14.575 2.805 ;
        RECT 14.865 2.635 15.035 2.805 ;
        RECT 15.325 2.635 15.495 2.805 ;
        RECT 15.785 2.635 15.955 2.805 ;
        RECT 16.245 2.635 16.415 2.805 ;
        RECT 16.705 2.635 16.875 2.805 ;
        RECT 17.165 2.635 17.335 2.805 ;
        RECT 17.625 2.635 17.795 2.805 ;
        RECT 18.085 2.635 18.255 2.805 ;
        RECT 18.545 2.635 18.715 2.805 ;
        RECT 19.005 2.635 19.175 2.805 ;
        RECT 19.465 2.635 19.635 2.805 ;
        RECT 19.925 2.635 20.095 2.805 ;
        RECT 20.385 2.635 20.555 2.805 ;
        RECT 20.845 2.635 21.015 2.805 ;
        RECT 21.305 2.635 21.475 2.805 ;
        RECT 21.765 2.635 21.935 2.805 ;
        RECT 22.225 2.635 22.395 2.805 ;
        RECT 22.685 2.635 22.855 2.805 ;
        RECT 23.145 2.635 23.315 2.805 ;
        RECT 23.605 2.635 23.775 2.805 ;
        RECT 24.065 2.635 24.235 2.805 ;
        RECT 24.525 2.635 24.695 2.805 ;
        RECT 24.985 2.635 25.155 2.805 ;
        RECT 25.445 2.635 25.615 2.805 ;
        RECT 1.525 1.785 1.695 1.955 ;
        RECT 4.745 1.785 4.915 1.955 ;
        RECT 7.965 1.785 8.135 1.955 ;
        RECT 11.185 1.785 11.355 1.955 ;
        RECT 14.405 1.785 14.575 1.955 ;
        RECT 17.625 1.785 17.795 1.955 ;
        RECT 20.845 1.785 21.015 1.955 ;
        RECT 24.065 1.785 24.235 1.955 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
        RECT 14.405 -0.085 14.575 0.085 ;
        RECT 14.865 -0.085 15.035 0.085 ;
        RECT 15.325 -0.085 15.495 0.085 ;
        RECT 15.785 -0.085 15.955 0.085 ;
        RECT 16.245 -0.085 16.415 0.085 ;
        RECT 16.705 -0.085 16.875 0.085 ;
        RECT 17.165 -0.085 17.335 0.085 ;
        RECT 17.625 -0.085 17.795 0.085 ;
        RECT 18.085 -0.085 18.255 0.085 ;
        RECT 18.545 -0.085 18.715 0.085 ;
        RECT 19.005 -0.085 19.175 0.085 ;
        RECT 19.465 -0.085 19.635 0.085 ;
        RECT 19.925 -0.085 20.095 0.085 ;
        RECT 20.385 -0.085 20.555 0.085 ;
        RECT 20.845 -0.085 21.015 0.085 ;
        RECT 21.305 -0.085 21.475 0.085 ;
        RECT 21.765 -0.085 21.935 0.085 ;
        RECT 22.225 -0.085 22.395 0.085 ;
        RECT 22.685 -0.085 22.855 0.085 ;
        RECT 23.145 -0.085 23.315 0.085 ;
        RECT 23.605 -0.085 23.775 0.085 ;
        RECT 24.065 -0.085 24.235 0.085 ;
        RECT 24.525 -0.085 24.695 0.085 ;
        RECT 24.985 -0.085 25.155 0.085 ;
        RECT 25.445 -0.085 25.615 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__muxb8to1_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__muxb8to1_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__muxb8to1_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.840 BY 5.440 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 18.795 4.115 20.185 4.385 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 18.795 1.055 20.185 1.325 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 17.075 4.115 18.465 4.385 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 17.075 1.055 18.465 1.325 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 6.375 4.115 7.765 4.385 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 6.375 1.055 7.765 1.325 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 4.655 4.115 6.045 4.385 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 4.655 1.055 6.045 1.325 ;
    END
  END D[0]
  PIN S[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.733200 ;
    PORT
      LAYER li1 ;
        RECT 24.160 4.115 24.755 4.445 ;
    END
  END S[7]
  PIN S[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.733200 ;
    PORT
      LAYER li1 ;
        RECT 24.160 0.995 24.755 1.325 ;
    END
  END S[6]
  PIN S[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.733200 ;
    PORT
      LAYER li1 ;
        RECT 12.505 4.115 13.100 4.445 ;
    END
  END S[5]
  PIN S[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.733200 ;
    PORT
      LAYER li1 ;
        RECT 12.505 0.995 13.100 1.325 ;
    END
  END S[4]
  PIN S[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.733200 ;
    PORT
      LAYER li1 ;
        RECT 11.740 4.115 12.335 4.445 ;
    END
  END S[3]
  PIN S[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.733200 ;
    PORT
      LAYER li1 ;
        RECT 11.740 0.995 12.335 1.325 ;
    END
  END S[2]
  PIN S[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.733200 ;
    PORT
      LAYER li1 ;
        RECT 0.085 4.115 0.680 4.445 ;
    END
  END S[1]
  PIN S[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.733200 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.680 1.325 ;
    END
  END S[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 24.840 0.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 5.200 24.840 5.680 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 5.355 0.315 5.525 ;
        RECT 0.180 5.335 0.315 5.355 ;
        RECT 6.125 5.335 6.295 5.525 ;
        RECT 18.545 5.335 18.715 5.525 ;
        RECT 0.180 5.240 1.530 5.335 ;
        RECT 4.095 5.240 8.325 5.335 ;
        RECT 10.890 5.240 13.950 5.335 ;
        RECT 16.515 5.240 20.745 5.335 ;
        RECT 23.310 5.240 24.660 5.335 ;
        RECT 0.180 4.655 24.660 5.240 ;
        RECT 1.895 4.460 10.525 4.655 ;
        RECT 14.315 4.460 22.945 4.655 ;
        RECT 4.095 4.425 8.325 4.460 ;
        RECT 16.515 4.425 20.745 4.460 ;
    END
    PORT
      LAYER pwell ;
        RECT 4.095 0.980 8.325 1.015 ;
        RECT 16.515 0.980 20.745 1.015 ;
        RECT 1.895 0.785 10.525 0.980 ;
        RECT 14.315 0.785 22.945 0.980 ;
        RECT 0.180 0.200 24.660 0.785 ;
        RECT 0.180 0.105 1.530 0.200 ;
        RECT 4.095 0.105 8.325 0.200 ;
        RECT 10.890 0.105 13.950 0.200 ;
        RECT 16.515 0.105 20.745 0.200 ;
        RECT 23.310 0.105 24.660 0.200 ;
        RECT 0.180 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 6.125 -0.085 6.295 0.105 ;
        RECT 18.545 -0.085 18.715 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 25.030 4.135 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 24.840 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.051200 ;
    PORT
      LAYER met1 ;
        RECT 2.225 3.640 2.515 3.685 ;
        RECT 3.165 3.640 3.455 3.685 ;
        RECT 8.965 3.640 9.255 3.685 ;
        RECT 9.905 3.640 10.195 3.685 ;
        RECT 14.645 3.640 14.935 3.685 ;
        RECT 15.585 3.640 15.875 3.685 ;
        RECT 21.385 3.640 21.675 3.685 ;
        RECT 22.325 3.640 22.615 3.685 ;
        RECT 2.225 3.500 22.615 3.640 ;
        RECT 2.225 3.455 2.515 3.500 ;
        RECT 3.165 3.455 3.455 3.500 ;
        RECT 8.965 3.455 9.255 3.500 ;
        RECT 9.905 3.455 10.195 3.500 ;
        RECT 14.645 3.455 14.935 3.500 ;
        RECT 15.585 3.455 15.875 3.500 ;
        RECT 21.385 3.455 21.675 3.500 ;
        RECT 22.325 3.455 22.615 3.500 ;
        RECT 2.225 1.940 2.515 1.985 ;
        RECT 3.165 1.940 3.455 1.985 ;
        RECT 8.965 1.940 9.255 1.985 ;
        RECT 9.905 1.940 10.195 1.985 ;
        RECT 14.645 1.940 14.935 1.985 ;
        RECT 15.585 1.940 15.875 1.985 ;
        RECT 21.385 1.940 21.675 1.985 ;
        RECT 22.325 1.940 22.615 1.985 ;
        RECT 2.225 1.800 22.615 1.940 ;
        RECT 2.225 1.755 2.515 1.800 ;
        RECT 3.165 1.755 3.455 1.800 ;
        RECT 8.965 1.755 9.255 1.800 ;
        RECT 9.905 1.755 10.195 1.800 ;
        RECT 14.645 1.755 14.935 1.800 ;
        RECT 15.585 1.755 15.875 1.800 ;
        RECT 21.385 1.755 21.675 1.800 ;
        RECT 22.325 1.755 22.615 1.800 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 5.355 24.840 5.525 ;
        RECT 0.270 4.830 0.560 5.355 ;
        RECT 0.770 4.615 1.020 5.160 ;
        RECT 1.190 4.830 1.480 5.355 ;
        RECT 1.985 5.015 4.015 5.185 ;
        RECT 1.985 4.670 2.235 5.015 ;
        RECT 0.850 4.375 1.020 4.615 ;
        RECT 2.405 4.375 2.735 4.845 ;
        RECT 2.905 4.670 3.075 5.015 ;
        RECT 3.245 4.555 3.575 4.845 ;
        RECT 3.745 4.725 4.015 5.015 ;
        RECT 4.185 4.895 4.435 5.355 ;
        RECT 4.605 4.725 4.935 5.185 ;
        RECT 5.105 4.895 5.375 5.355 ;
        RECT 5.545 4.725 5.875 5.185 ;
        RECT 3.745 4.555 5.875 4.725 ;
        RECT 6.045 4.555 6.375 5.355 ;
        RECT 6.545 4.725 6.875 5.185 ;
        RECT 7.045 4.895 7.315 5.355 ;
        RECT 7.485 4.725 7.815 5.185 ;
        RECT 7.985 4.895 8.235 5.355 ;
        RECT 8.405 5.015 10.435 5.185 ;
        RECT 8.405 4.725 8.675 5.015 ;
        RECT 6.545 4.555 8.675 4.725 ;
        RECT 8.845 4.555 9.175 4.845 ;
        RECT 9.345 4.670 9.515 5.015 ;
        RECT 3.245 4.375 3.475 4.555 ;
        RECT 0.850 4.045 2.035 4.375 ;
        RECT 2.205 4.075 3.475 4.375 ;
        RECT 0.850 3.835 1.020 4.045 ;
        RECT 0.220 2.805 0.520 3.835 ;
        RECT 0.690 2.975 1.020 3.835 ;
        RECT 1.215 2.805 1.490 3.835 ;
        RECT 1.735 2.975 2.035 3.875 ;
        RECT 0.000 2.635 2.035 2.805 ;
        RECT 0.220 1.605 0.520 2.635 ;
        RECT 0.690 1.605 1.020 2.465 ;
        RECT 1.215 1.605 1.490 2.635 ;
        RECT 0.850 1.395 1.020 1.605 ;
        RECT 1.735 1.565 2.035 2.465 ;
        RECT 0.850 1.065 2.035 1.395 ;
        RECT 2.205 1.365 2.535 4.075 ;
        RECT 2.705 2.975 2.975 3.905 ;
        RECT 2.705 1.535 2.975 2.465 ;
        RECT 3.145 1.365 3.475 4.075 ;
        RECT 8.945 4.375 9.175 4.555 ;
        RECT 9.685 4.375 10.015 4.845 ;
        RECT 10.185 4.670 10.435 5.015 ;
        RECT 10.940 4.830 11.230 5.355 ;
        RECT 11.400 4.615 11.650 5.160 ;
        RECT 11.860 4.830 12.150 5.355 ;
        RECT 12.690 4.830 12.980 5.355 ;
        RECT 13.190 4.615 13.440 5.160 ;
        RECT 13.610 4.830 13.900 5.355 ;
        RECT 14.405 5.015 16.435 5.185 ;
        RECT 14.405 4.670 14.655 5.015 ;
        RECT 11.400 4.375 11.570 4.615 ;
        RECT 8.945 4.075 10.215 4.375 ;
        RECT 3.645 3.775 5.875 3.945 ;
        RECT 3.645 2.975 3.945 3.775 ;
        RECT 4.165 2.805 4.435 3.605 ;
        RECT 4.605 2.975 4.935 3.775 ;
        RECT 5.105 2.805 5.375 3.605 ;
        RECT 5.545 2.975 5.875 3.775 ;
        RECT 6.045 2.805 6.375 3.945 ;
        RECT 6.545 3.775 8.775 3.945 ;
        RECT 6.545 2.975 6.875 3.775 ;
        RECT 7.045 2.805 7.315 3.605 ;
        RECT 7.485 2.975 7.815 3.775 ;
        RECT 7.985 2.805 8.255 3.605 ;
        RECT 8.475 2.975 8.775 3.775 ;
        RECT 3.645 2.635 8.775 2.805 ;
        RECT 3.645 1.665 3.945 2.465 ;
        RECT 4.165 1.835 4.435 2.635 ;
        RECT 4.605 1.665 4.935 2.465 ;
        RECT 5.105 1.835 5.375 2.635 ;
        RECT 5.545 1.665 5.875 2.465 ;
        RECT 3.645 1.495 5.875 1.665 ;
        RECT 6.045 1.495 6.375 2.635 ;
        RECT 6.545 1.665 6.875 2.465 ;
        RECT 7.045 1.835 7.315 2.635 ;
        RECT 7.485 1.665 7.815 2.465 ;
        RECT 7.985 1.835 8.255 2.635 ;
        RECT 8.475 1.665 8.775 2.465 ;
        RECT 6.545 1.495 8.775 1.665 ;
        RECT 2.205 1.065 3.475 1.365 ;
        RECT 0.850 0.825 1.020 1.065 ;
        RECT 0.270 0.085 0.560 0.610 ;
        RECT 0.770 0.280 1.020 0.825 ;
        RECT 1.190 0.085 1.480 0.610 ;
        RECT 1.985 0.425 2.235 0.770 ;
        RECT 2.405 0.595 2.735 1.065 ;
        RECT 3.245 0.885 3.475 1.065 ;
        RECT 8.945 1.365 9.275 4.075 ;
        RECT 9.445 2.975 9.715 3.905 ;
        RECT 9.445 1.535 9.715 2.465 ;
        RECT 9.885 1.365 10.215 4.075 ;
        RECT 10.385 4.045 11.570 4.375 ;
        RECT 10.385 2.975 10.685 3.875 ;
        RECT 11.400 3.835 11.570 4.045 ;
        RECT 13.270 4.375 13.440 4.615 ;
        RECT 14.825 4.375 15.155 4.845 ;
        RECT 15.325 4.670 15.495 5.015 ;
        RECT 15.665 4.555 15.995 4.845 ;
        RECT 16.165 4.725 16.435 5.015 ;
        RECT 16.605 4.895 16.855 5.355 ;
        RECT 17.025 4.725 17.355 5.185 ;
        RECT 17.525 4.895 17.795 5.355 ;
        RECT 17.965 4.725 18.295 5.185 ;
        RECT 16.165 4.555 18.295 4.725 ;
        RECT 18.465 4.555 18.795 5.355 ;
        RECT 18.965 4.725 19.295 5.185 ;
        RECT 19.465 4.895 19.735 5.355 ;
        RECT 19.905 4.725 20.235 5.185 ;
        RECT 20.405 4.895 20.655 5.355 ;
        RECT 20.825 5.015 22.855 5.185 ;
        RECT 20.825 4.725 21.095 5.015 ;
        RECT 18.965 4.555 21.095 4.725 ;
        RECT 21.265 4.555 21.595 4.845 ;
        RECT 21.765 4.670 21.935 5.015 ;
        RECT 15.665 4.375 15.895 4.555 ;
        RECT 13.270 4.045 14.455 4.375 ;
        RECT 14.625 4.075 15.895 4.375 ;
        RECT 13.270 3.835 13.440 4.045 ;
        RECT 10.930 2.805 11.205 3.835 ;
        RECT 11.400 2.975 11.730 3.835 ;
        RECT 11.900 2.805 12.200 3.835 ;
        RECT 12.640 2.805 12.940 3.835 ;
        RECT 13.110 2.975 13.440 3.835 ;
        RECT 13.635 2.805 13.910 3.835 ;
        RECT 14.155 2.975 14.455 3.875 ;
        RECT 10.385 2.635 14.455 2.805 ;
        RECT 10.385 1.565 10.685 2.465 ;
        RECT 10.930 1.605 11.205 2.635 ;
        RECT 11.400 1.605 11.730 2.465 ;
        RECT 11.900 1.605 12.200 2.635 ;
        RECT 12.640 1.605 12.940 2.635 ;
        RECT 13.110 1.605 13.440 2.465 ;
        RECT 13.635 1.605 13.910 2.635 ;
        RECT 11.400 1.395 11.570 1.605 ;
        RECT 8.945 1.065 10.215 1.365 ;
        RECT 10.385 1.065 11.570 1.395 ;
        RECT 8.945 0.885 9.175 1.065 ;
        RECT 2.905 0.425 3.075 0.770 ;
        RECT 3.245 0.595 3.575 0.885 ;
        RECT 3.745 0.715 5.875 0.885 ;
        RECT 3.745 0.425 4.015 0.715 ;
        RECT 1.985 0.255 4.015 0.425 ;
        RECT 4.185 0.085 4.435 0.545 ;
        RECT 4.605 0.255 4.935 0.715 ;
        RECT 5.105 0.085 5.375 0.545 ;
        RECT 5.545 0.255 5.875 0.715 ;
        RECT 6.045 0.085 6.375 0.885 ;
        RECT 6.545 0.715 8.675 0.885 ;
        RECT 6.545 0.255 6.875 0.715 ;
        RECT 7.045 0.085 7.315 0.545 ;
        RECT 7.485 0.255 7.815 0.715 ;
        RECT 7.985 0.085 8.235 0.545 ;
        RECT 8.405 0.425 8.675 0.715 ;
        RECT 8.845 0.595 9.175 0.885 ;
        RECT 9.345 0.425 9.515 0.770 ;
        RECT 9.685 0.595 10.015 1.065 ;
        RECT 11.400 0.825 11.570 1.065 ;
        RECT 13.270 1.395 13.440 1.605 ;
        RECT 14.155 1.565 14.455 2.465 ;
        RECT 13.270 1.065 14.455 1.395 ;
        RECT 14.625 1.365 14.955 4.075 ;
        RECT 15.125 2.975 15.395 3.905 ;
        RECT 15.125 1.535 15.395 2.465 ;
        RECT 15.565 1.365 15.895 4.075 ;
        RECT 21.365 4.375 21.595 4.555 ;
        RECT 22.105 4.375 22.435 4.845 ;
        RECT 22.605 4.670 22.855 5.015 ;
        RECT 23.360 4.830 23.650 5.355 ;
        RECT 23.820 4.615 24.070 5.160 ;
        RECT 24.280 4.830 24.570 5.355 ;
        RECT 23.820 4.375 23.990 4.615 ;
        RECT 21.365 4.075 22.635 4.375 ;
        RECT 16.065 3.775 18.295 3.945 ;
        RECT 16.065 2.975 16.365 3.775 ;
        RECT 16.585 2.805 16.855 3.605 ;
        RECT 17.025 2.975 17.355 3.775 ;
        RECT 17.525 2.805 17.795 3.605 ;
        RECT 17.965 2.975 18.295 3.775 ;
        RECT 18.465 2.805 18.795 3.945 ;
        RECT 18.965 3.775 21.195 3.945 ;
        RECT 18.965 2.975 19.295 3.775 ;
        RECT 19.465 2.805 19.735 3.605 ;
        RECT 19.905 2.975 20.235 3.775 ;
        RECT 20.405 2.805 20.675 3.605 ;
        RECT 20.895 2.975 21.195 3.775 ;
        RECT 16.065 2.635 21.195 2.805 ;
        RECT 16.065 1.665 16.365 2.465 ;
        RECT 16.585 1.835 16.855 2.635 ;
        RECT 17.025 1.665 17.355 2.465 ;
        RECT 17.525 1.835 17.795 2.635 ;
        RECT 17.965 1.665 18.295 2.465 ;
        RECT 16.065 1.495 18.295 1.665 ;
        RECT 18.465 1.495 18.795 2.635 ;
        RECT 18.965 1.665 19.295 2.465 ;
        RECT 19.465 1.835 19.735 2.635 ;
        RECT 19.905 1.665 20.235 2.465 ;
        RECT 20.405 1.835 20.675 2.635 ;
        RECT 20.895 1.665 21.195 2.465 ;
        RECT 18.965 1.495 21.195 1.665 ;
        RECT 14.625 1.065 15.895 1.365 ;
        RECT 13.270 0.825 13.440 1.065 ;
        RECT 10.185 0.425 10.435 0.770 ;
        RECT 8.405 0.255 10.435 0.425 ;
        RECT 10.940 0.085 11.230 0.610 ;
        RECT 11.400 0.280 11.650 0.825 ;
        RECT 11.860 0.085 12.150 0.610 ;
        RECT 12.690 0.085 12.980 0.610 ;
        RECT 13.190 0.280 13.440 0.825 ;
        RECT 13.610 0.085 13.900 0.610 ;
        RECT 14.405 0.425 14.655 0.770 ;
        RECT 14.825 0.595 15.155 1.065 ;
        RECT 15.665 0.885 15.895 1.065 ;
        RECT 21.365 1.365 21.695 4.075 ;
        RECT 21.865 2.975 22.135 3.905 ;
        RECT 21.865 1.535 22.135 2.465 ;
        RECT 22.305 1.365 22.635 4.075 ;
        RECT 22.805 4.045 23.990 4.375 ;
        RECT 22.805 2.975 23.105 3.875 ;
        RECT 23.820 3.835 23.990 4.045 ;
        RECT 23.350 2.805 23.625 3.835 ;
        RECT 23.820 2.975 24.150 3.835 ;
        RECT 24.320 2.805 24.620 3.835 ;
        RECT 22.805 2.635 24.840 2.805 ;
        RECT 22.805 1.565 23.105 2.465 ;
        RECT 23.350 1.605 23.625 2.635 ;
        RECT 23.820 1.605 24.150 2.465 ;
        RECT 24.320 1.605 24.620 2.635 ;
        RECT 23.820 1.395 23.990 1.605 ;
        RECT 21.365 1.065 22.635 1.365 ;
        RECT 22.805 1.065 23.990 1.395 ;
        RECT 21.365 0.885 21.595 1.065 ;
        RECT 15.325 0.425 15.495 0.770 ;
        RECT 15.665 0.595 15.995 0.885 ;
        RECT 16.165 0.715 18.295 0.885 ;
        RECT 16.165 0.425 16.435 0.715 ;
        RECT 14.405 0.255 16.435 0.425 ;
        RECT 16.605 0.085 16.855 0.545 ;
        RECT 17.025 0.255 17.355 0.715 ;
        RECT 17.525 0.085 17.795 0.545 ;
        RECT 17.965 0.255 18.295 0.715 ;
        RECT 18.465 0.085 18.795 0.885 ;
        RECT 18.965 0.715 21.095 0.885 ;
        RECT 18.965 0.255 19.295 0.715 ;
        RECT 19.465 0.085 19.735 0.545 ;
        RECT 19.905 0.255 20.235 0.715 ;
        RECT 20.405 0.085 20.655 0.545 ;
        RECT 20.825 0.425 21.095 0.715 ;
        RECT 21.265 0.595 21.595 0.885 ;
        RECT 21.765 0.425 21.935 0.770 ;
        RECT 22.105 0.595 22.435 1.065 ;
        RECT 23.820 0.825 23.990 1.065 ;
        RECT 22.605 0.425 22.855 0.770 ;
        RECT 20.825 0.255 22.855 0.425 ;
        RECT 23.360 0.085 23.650 0.610 ;
        RECT 23.820 0.280 24.070 0.825 ;
        RECT 24.280 0.085 24.570 0.610 ;
        RECT 0.000 -0.085 24.840 0.085 ;
      LAYER mcon ;
        RECT 0.145 5.355 0.315 5.525 ;
        RECT 0.605 5.355 0.775 5.525 ;
        RECT 1.065 5.355 1.235 5.525 ;
        RECT 1.525 5.355 1.695 5.525 ;
        RECT 1.985 5.355 2.155 5.525 ;
        RECT 2.445 5.355 2.615 5.525 ;
        RECT 2.905 5.355 3.075 5.525 ;
        RECT 3.365 5.355 3.535 5.525 ;
        RECT 3.825 5.355 3.995 5.525 ;
        RECT 4.285 5.355 4.455 5.525 ;
        RECT 4.745 5.355 4.915 5.525 ;
        RECT 5.205 5.355 5.375 5.525 ;
        RECT 5.665 5.355 5.835 5.525 ;
        RECT 6.125 5.355 6.295 5.525 ;
        RECT 6.585 5.355 6.755 5.525 ;
        RECT 7.045 5.355 7.215 5.525 ;
        RECT 7.505 5.355 7.675 5.525 ;
        RECT 7.965 5.355 8.135 5.525 ;
        RECT 8.425 5.355 8.595 5.525 ;
        RECT 8.885 5.355 9.055 5.525 ;
        RECT 9.345 5.355 9.515 5.525 ;
        RECT 9.805 5.355 9.975 5.525 ;
        RECT 10.265 5.355 10.435 5.525 ;
        RECT 10.725 5.355 10.895 5.525 ;
        RECT 11.185 5.355 11.355 5.525 ;
        RECT 11.645 5.355 11.815 5.525 ;
        RECT 12.105 5.355 12.275 5.525 ;
        RECT 12.565 5.355 12.735 5.525 ;
        RECT 13.025 5.355 13.195 5.525 ;
        RECT 13.485 5.355 13.655 5.525 ;
        RECT 13.945 5.355 14.115 5.525 ;
        RECT 14.405 5.355 14.575 5.525 ;
        RECT 14.865 5.355 15.035 5.525 ;
        RECT 15.325 5.355 15.495 5.525 ;
        RECT 15.785 5.355 15.955 5.525 ;
        RECT 16.245 5.355 16.415 5.525 ;
        RECT 16.705 5.355 16.875 5.525 ;
        RECT 17.165 5.355 17.335 5.525 ;
        RECT 17.625 5.355 17.795 5.525 ;
        RECT 18.085 5.355 18.255 5.525 ;
        RECT 18.545 5.355 18.715 5.525 ;
        RECT 19.005 5.355 19.175 5.525 ;
        RECT 19.465 5.355 19.635 5.525 ;
        RECT 19.925 5.355 20.095 5.525 ;
        RECT 20.385 5.355 20.555 5.525 ;
        RECT 20.845 5.355 21.015 5.525 ;
        RECT 21.305 5.355 21.475 5.525 ;
        RECT 21.765 5.355 21.935 5.525 ;
        RECT 22.225 5.355 22.395 5.525 ;
        RECT 22.685 5.355 22.855 5.525 ;
        RECT 23.145 5.355 23.315 5.525 ;
        RECT 23.605 5.355 23.775 5.525 ;
        RECT 24.065 5.355 24.235 5.525 ;
        RECT 24.525 5.355 24.695 5.525 ;
        RECT 1.805 3.130 1.975 3.300 ;
        RECT 2.285 3.485 2.455 3.655 ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.805 2.140 1.975 2.310 ;
        RECT 2.755 3.130 2.925 3.300 ;
        RECT 3.225 3.485 3.395 3.655 ;
        RECT 2.285 1.785 2.455 1.955 ;
        RECT 2.755 2.140 2.925 2.310 ;
        RECT 3.705 3.130 3.875 3.300 ;
        RECT 4.685 3.130 4.855 3.300 ;
        RECT 5.625 3.130 5.795 3.300 ;
        RECT 6.625 3.130 6.795 3.300 ;
        RECT 7.565 3.130 7.735 3.300 ;
        RECT 8.545 3.130 8.715 3.300 ;
        RECT 9.025 3.485 9.195 3.655 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 3.225 1.785 3.395 1.955 ;
        RECT 3.705 2.140 3.875 2.310 ;
        RECT 4.685 2.140 4.855 2.310 ;
        RECT 5.625 2.140 5.795 2.310 ;
        RECT 6.625 2.140 6.795 2.310 ;
        RECT 7.565 2.140 7.735 2.310 ;
        RECT 8.545 2.140 8.715 2.310 ;
        RECT 9.495 3.130 9.665 3.300 ;
        RECT 9.965 3.485 10.135 3.655 ;
        RECT 9.025 1.785 9.195 1.955 ;
        RECT 9.495 2.140 9.665 2.310 ;
        RECT 10.445 3.130 10.615 3.300 ;
        RECT 14.225 3.130 14.395 3.300 ;
        RECT 14.705 3.485 14.875 3.655 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 9.965 1.785 10.135 1.955 ;
        RECT 10.445 2.140 10.615 2.310 ;
        RECT 14.225 2.140 14.395 2.310 ;
        RECT 15.175 3.130 15.345 3.300 ;
        RECT 15.645 3.485 15.815 3.655 ;
        RECT 14.705 1.785 14.875 1.955 ;
        RECT 15.175 2.140 15.345 2.310 ;
        RECT 16.125 3.130 16.295 3.300 ;
        RECT 17.105 3.130 17.275 3.300 ;
        RECT 18.045 3.130 18.215 3.300 ;
        RECT 19.045 3.130 19.215 3.300 ;
        RECT 19.985 3.130 20.155 3.300 ;
        RECT 20.965 3.130 21.135 3.300 ;
        RECT 21.445 3.485 21.615 3.655 ;
        RECT 16.245 2.635 16.415 2.805 ;
        RECT 16.705 2.635 16.875 2.805 ;
        RECT 17.165 2.635 17.335 2.805 ;
        RECT 17.625 2.635 17.795 2.805 ;
        RECT 18.085 2.635 18.255 2.805 ;
        RECT 18.545 2.635 18.715 2.805 ;
        RECT 19.005 2.635 19.175 2.805 ;
        RECT 19.465 2.635 19.635 2.805 ;
        RECT 19.925 2.635 20.095 2.805 ;
        RECT 20.385 2.635 20.555 2.805 ;
        RECT 20.845 2.635 21.015 2.805 ;
        RECT 15.645 1.785 15.815 1.955 ;
        RECT 16.125 2.140 16.295 2.310 ;
        RECT 17.105 2.140 17.275 2.310 ;
        RECT 18.045 2.140 18.215 2.310 ;
        RECT 19.045 2.140 19.215 2.310 ;
        RECT 19.985 2.140 20.155 2.310 ;
        RECT 20.965 2.140 21.135 2.310 ;
        RECT 21.915 3.130 22.085 3.300 ;
        RECT 22.385 3.485 22.555 3.655 ;
        RECT 21.445 1.785 21.615 1.955 ;
        RECT 21.915 2.140 22.085 2.310 ;
        RECT 22.865 3.130 23.035 3.300 ;
        RECT 23.145 2.635 23.315 2.805 ;
        RECT 23.605 2.635 23.775 2.805 ;
        RECT 24.065 2.635 24.235 2.805 ;
        RECT 24.525 2.635 24.695 2.805 ;
        RECT 22.385 1.785 22.555 1.955 ;
        RECT 22.865 2.140 23.035 2.310 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
        RECT 14.405 -0.085 14.575 0.085 ;
        RECT 14.865 -0.085 15.035 0.085 ;
        RECT 15.325 -0.085 15.495 0.085 ;
        RECT 15.785 -0.085 15.955 0.085 ;
        RECT 16.245 -0.085 16.415 0.085 ;
        RECT 16.705 -0.085 16.875 0.085 ;
        RECT 17.165 -0.085 17.335 0.085 ;
        RECT 17.625 -0.085 17.795 0.085 ;
        RECT 18.085 -0.085 18.255 0.085 ;
        RECT 18.545 -0.085 18.715 0.085 ;
        RECT 19.005 -0.085 19.175 0.085 ;
        RECT 19.465 -0.085 19.635 0.085 ;
        RECT 19.925 -0.085 20.095 0.085 ;
        RECT 20.385 -0.085 20.555 0.085 ;
        RECT 20.845 -0.085 21.015 0.085 ;
        RECT 21.305 -0.085 21.475 0.085 ;
        RECT 21.765 -0.085 21.935 0.085 ;
        RECT 22.225 -0.085 22.395 0.085 ;
        RECT 22.685 -0.085 22.855 0.085 ;
        RECT 23.145 -0.085 23.315 0.085 ;
        RECT 23.605 -0.085 23.775 0.085 ;
        RECT 24.065 -0.085 24.235 0.085 ;
        RECT 24.525 -0.085 24.695 0.085 ;
      LAYER met1 ;
        RECT 1.745 3.285 2.035 3.330 ;
        RECT 2.695 3.285 2.985 3.330 ;
        RECT 3.645 3.285 3.935 3.330 ;
        RECT 4.625 3.285 4.915 3.330 ;
        RECT 5.565 3.285 5.855 3.330 ;
        RECT 1.745 3.145 5.855 3.285 ;
        RECT 1.745 3.100 2.035 3.145 ;
        RECT 2.695 3.100 2.985 3.145 ;
        RECT 3.645 3.100 3.935 3.145 ;
        RECT 4.625 3.100 4.915 3.145 ;
        RECT 5.565 3.100 5.855 3.145 ;
        RECT 6.565 3.285 6.855 3.330 ;
        RECT 7.505 3.285 7.795 3.330 ;
        RECT 8.485 3.285 8.775 3.330 ;
        RECT 9.435 3.285 9.725 3.330 ;
        RECT 10.385 3.285 10.675 3.330 ;
        RECT 6.565 3.145 10.675 3.285 ;
        RECT 6.565 3.100 6.855 3.145 ;
        RECT 7.505 3.100 7.795 3.145 ;
        RECT 8.485 3.100 8.775 3.145 ;
        RECT 9.435 3.100 9.725 3.145 ;
        RECT 10.385 3.100 10.675 3.145 ;
        RECT 14.165 3.285 14.455 3.330 ;
        RECT 15.115 3.285 15.405 3.330 ;
        RECT 16.065 3.285 16.355 3.330 ;
        RECT 17.045 3.285 17.335 3.330 ;
        RECT 17.985 3.285 18.275 3.330 ;
        RECT 14.165 3.145 18.275 3.285 ;
        RECT 14.165 3.100 14.455 3.145 ;
        RECT 15.115 3.100 15.405 3.145 ;
        RECT 16.065 3.100 16.355 3.145 ;
        RECT 17.045 3.100 17.335 3.145 ;
        RECT 17.985 3.100 18.275 3.145 ;
        RECT 18.985 3.285 19.275 3.330 ;
        RECT 19.925 3.285 20.215 3.330 ;
        RECT 20.905 3.285 21.195 3.330 ;
        RECT 21.855 3.285 22.145 3.330 ;
        RECT 22.805 3.285 23.095 3.330 ;
        RECT 18.985 3.145 23.095 3.285 ;
        RECT 18.985 3.100 19.275 3.145 ;
        RECT 19.925 3.100 20.215 3.145 ;
        RECT 20.905 3.100 21.195 3.145 ;
        RECT 21.855 3.100 22.145 3.145 ;
        RECT 22.805 3.100 23.095 3.145 ;
        RECT 1.745 2.295 2.035 2.340 ;
        RECT 2.695 2.295 2.985 2.340 ;
        RECT 3.645 2.295 3.935 2.340 ;
        RECT 4.625 2.295 4.915 2.340 ;
        RECT 5.565 2.295 5.855 2.340 ;
        RECT 1.745 2.155 5.855 2.295 ;
        RECT 1.745 2.110 2.035 2.155 ;
        RECT 2.695 2.110 2.985 2.155 ;
        RECT 3.645 2.110 3.935 2.155 ;
        RECT 4.625 2.110 4.915 2.155 ;
        RECT 5.565 2.110 5.855 2.155 ;
        RECT 6.565 2.295 6.855 2.340 ;
        RECT 7.505 2.295 7.795 2.340 ;
        RECT 8.485 2.295 8.775 2.340 ;
        RECT 9.435 2.295 9.725 2.340 ;
        RECT 10.385 2.295 10.675 2.340 ;
        RECT 6.565 2.155 10.675 2.295 ;
        RECT 6.565 2.110 6.855 2.155 ;
        RECT 7.505 2.110 7.795 2.155 ;
        RECT 8.485 2.110 8.775 2.155 ;
        RECT 9.435 2.110 9.725 2.155 ;
        RECT 10.385 2.110 10.675 2.155 ;
        RECT 14.165 2.295 14.455 2.340 ;
        RECT 15.115 2.295 15.405 2.340 ;
        RECT 16.065 2.295 16.355 2.340 ;
        RECT 17.045 2.295 17.335 2.340 ;
        RECT 17.985 2.295 18.275 2.340 ;
        RECT 14.165 2.155 18.275 2.295 ;
        RECT 14.165 2.110 14.455 2.155 ;
        RECT 15.115 2.110 15.405 2.155 ;
        RECT 16.065 2.110 16.355 2.155 ;
        RECT 17.045 2.110 17.335 2.155 ;
        RECT 17.985 2.110 18.275 2.155 ;
        RECT 18.985 2.295 19.275 2.340 ;
        RECT 19.925 2.295 20.215 2.340 ;
        RECT 20.905 2.295 21.195 2.340 ;
        RECT 21.855 2.295 22.145 2.340 ;
        RECT 22.805 2.295 23.095 2.340 ;
        RECT 18.985 2.155 23.095 2.295 ;
        RECT 18.985 2.110 19.275 2.155 ;
        RECT 19.925 2.110 20.215 2.155 ;
        RECT 20.905 2.110 21.195 2.155 ;
        RECT 21.855 2.110 22.145 2.155 ;
        RECT 22.805 2.110 23.095 2.155 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__muxb8to1_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__muxb16to1_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__muxb16to1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.020 BY 5.440 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 16.185 4.815 16.460 5.045 ;
        RECT 16.290 4.385 16.460 4.815 ;
        RECT 16.290 4.115 16.685 4.385 ;
    END
  END D[15]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 12.980 4.815 13.255 5.045 ;
        RECT 12.980 4.385 13.150 4.815 ;
        RECT 12.755 4.115 13.150 4.385 ;
    END
  END D[14]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 12.045 4.815 12.320 5.045 ;
        RECT 12.150 4.385 12.320 4.815 ;
        RECT 12.150 4.115 12.545 4.385 ;
    END
  END D[13]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 8.840 4.815 9.115 5.045 ;
        RECT 8.840 4.385 9.010 4.815 ;
        RECT 8.615 4.115 9.010 4.385 ;
    END
  END D[12]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 7.905 4.815 8.180 5.045 ;
        RECT 8.010 4.385 8.180 4.815 ;
        RECT 8.010 4.115 8.405 4.385 ;
    END
  END D[11]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 4.700 4.815 4.975 5.045 ;
        RECT 4.700 4.385 4.870 4.815 ;
        RECT 4.475 4.115 4.870 4.385 ;
    END
  END D[10]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 3.765 4.815 4.040 5.045 ;
        RECT 3.870 4.385 4.040 4.815 ;
        RECT 3.870 4.115 4.265 4.385 ;
    END
  END D[9]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.560 4.815 0.835 5.045 ;
        RECT 0.560 4.385 0.730 4.815 ;
        RECT 0.335 4.115 0.730 4.385 ;
    END
  END D[8]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 16.290 1.055 16.685 1.325 ;
        RECT 16.290 0.625 16.460 1.055 ;
        RECT 16.185 0.395 16.460 0.625 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 12.755 1.055 13.150 1.325 ;
        RECT 12.980 0.625 13.150 1.055 ;
        RECT 12.980 0.395 13.255 0.625 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 12.150 1.055 12.545 1.325 ;
        RECT 12.150 0.625 12.320 1.055 ;
        RECT 12.045 0.395 12.320 0.625 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 8.615 1.055 9.010 1.325 ;
        RECT 8.840 0.625 9.010 1.055 ;
        RECT 8.840 0.395 9.115 0.625 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 8.010 1.055 8.405 1.325 ;
        RECT 8.010 0.625 8.180 1.055 ;
        RECT 7.905 0.395 8.180 0.625 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 4.475 1.055 4.870 1.325 ;
        RECT 4.700 0.625 4.870 1.055 ;
        RECT 4.700 0.395 4.975 0.625 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 3.870 1.055 4.265 1.325 ;
        RECT 3.870 0.625 4.040 1.055 ;
        RECT 3.765 0.395 4.040 0.625 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.335 1.055 0.730 1.325 ;
        RECT 0.560 0.625 0.730 1.055 ;
        RECT 0.560 0.395 0.835 0.625 ;
    END
  END D[0]
  PIN S[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 14.815 4.145 15.215 4.495 ;
    END
  END S[15]
  PIN S[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 14.225 4.145 14.625 4.495 ;
    END
  END S[14]
  PIN S[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 10.675 4.145 11.075 4.495 ;
    END
  END S[13]
  PIN S[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 10.085 4.145 10.485 4.495 ;
    END
  END S[12]
  PIN S[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 6.535 4.145 6.935 4.495 ;
    END
  END S[11]
  PIN S[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 5.945 4.145 6.345 4.495 ;
    END
  END S[10]
  PIN S[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 2.395 4.145 2.795 4.495 ;
    END
  END S[9]
  PIN S[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 1.805 4.145 2.205 4.495 ;
    END
  END S[8]
  PIN S[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 14.815 0.945 15.215 1.295 ;
    END
  END S[7]
  PIN S[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 14.225 0.945 14.625 1.295 ;
    END
  END S[6]
  PIN S[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 10.675 0.945 11.075 1.295 ;
    END
  END S[5]
  PIN S[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 10.085 0.945 10.485 1.295 ;
    END
  END S[4]
  PIN S[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 6.535 0.945 6.935 1.295 ;
    END
  END S[3]
  PIN S[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 5.945 0.945 6.345 1.295 ;
    END
  END S[2]
  PIN S[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 2.395 0.945 2.795 1.295 ;
    END
  END S[1]
  PIN S[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 1.805 0.945 2.205 1.295 ;
    END
  END S[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 17.020 0.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 5.200 17.020 5.680 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 5.335 0.315 5.525 ;
        RECT 4.285 5.335 4.455 5.525 ;
        RECT 8.425 5.335 8.595 5.525 ;
        RECT 12.565 5.335 12.735 5.525 ;
        RECT 16.705 5.335 16.875 5.525 ;
        RECT 0.005 4.555 17.015 5.335 ;
        RECT 0.005 4.425 0.925 4.555 ;
        RECT 3.675 4.425 5.065 4.555 ;
        RECT 7.815 4.425 9.205 4.555 ;
        RECT 11.955 4.425 13.345 4.555 ;
        RECT 16.095 4.425 17.015 4.555 ;
    END
    PORT
      LAYER pwell ;
        RECT 0.005 0.885 0.925 1.015 ;
        RECT 3.675 0.885 5.065 1.015 ;
        RECT 7.815 0.885 9.205 1.015 ;
        RECT 11.955 0.885 13.345 1.015 ;
        RECT 16.095 0.885 17.015 1.015 ;
        RECT 0.005 0.105 17.015 0.885 ;
        RECT 0.145 -0.085 0.315 0.105 ;
        RECT 4.285 -0.085 4.455 0.105 ;
        RECT 8.425 -0.085 8.595 0.105 ;
        RECT 12.565 -0.085 12.735 0.105 ;
        RECT 16.705 -0.085 16.875 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 17.210 4.135 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 17.020 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.705600 ;
    PORT
      LAYER met1 ;
        RECT 1.005 3.640 1.295 3.685 ;
        RECT 3.305 3.640 3.595 3.685 ;
        RECT 5.145 3.640 5.435 3.685 ;
        RECT 7.445 3.640 7.735 3.685 ;
        RECT 9.285 3.640 9.575 3.685 ;
        RECT 11.585 3.640 11.875 3.685 ;
        RECT 13.425 3.640 13.715 3.685 ;
        RECT 15.725 3.640 16.015 3.685 ;
        RECT 1.005 3.500 16.015 3.640 ;
        RECT 1.005 3.455 1.295 3.500 ;
        RECT 3.305 3.455 3.595 3.500 ;
        RECT 5.145 3.455 5.435 3.500 ;
        RECT 7.445 3.455 7.735 3.500 ;
        RECT 9.285 3.455 9.575 3.500 ;
        RECT 11.585 3.455 11.875 3.500 ;
        RECT 13.425 3.455 13.715 3.500 ;
        RECT 15.725 3.455 16.015 3.500 ;
        RECT 1.005 1.940 1.295 1.985 ;
        RECT 3.305 1.940 3.595 1.985 ;
        RECT 5.145 1.940 5.435 1.985 ;
        RECT 7.445 1.940 7.735 1.985 ;
        RECT 9.285 1.940 9.575 1.985 ;
        RECT 11.585 1.940 11.875 1.985 ;
        RECT 13.425 1.940 13.715 1.985 ;
        RECT 15.725 1.940 16.015 1.985 ;
        RECT 1.005 1.800 16.015 1.940 ;
        RECT 1.005 1.755 1.295 1.800 ;
        RECT 3.305 1.755 3.595 1.800 ;
        RECT 5.145 1.755 5.435 1.800 ;
        RECT 7.445 1.755 7.735 1.800 ;
        RECT 9.285 1.755 9.575 1.800 ;
        RECT 11.585 1.755 11.875 1.800 ;
        RECT 13.425 1.755 13.715 1.800 ;
        RECT 15.725 1.755 16.015 1.800 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 5.355 17.020 5.525 ;
        RECT 0.130 4.555 0.390 5.355 ;
        RECT 1.045 4.605 1.290 5.110 ;
        RECT 1.650 4.855 1.900 5.110 ;
        RECT 0.900 4.435 1.290 4.605 ;
        RECT 1.460 4.685 1.900 4.855 ;
        RECT 2.135 4.780 2.465 5.355 ;
        RECT 2.700 4.855 2.950 5.110 ;
        RECT 2.700 4.685 3.140 4.855 ;
        RECT 0.095 2.805 0.425 3.945 ;
        RECT 0.900 3.685 1.070 4.435 ;
        RECT 1.460 4.265 1.630 4.685 ;
        RECT 1.240 3.975 1.630 4.265 ;
        RECT 2.970 4.265 3.140 4.685 ;
        RECT 3.310 4.605 3.555 5.110 ;
        RECT 3.310 4.435 3.700 4.605 ;
        RECT 4.210 4.555 4.530 5.355 ;
        RECT 5.185 4.605 5.430 5.110 ;
        RECT 5.790 4.855 6.040 5.110 ;
        RECT 2.970 3.975 3.360 4.265 ;
        RECT 1.240 3.935 1.940 3.975 ;
        RECT 1.460 3.805 1.940 3.935 ;
        RECT 0.900 3.635 1.295 3.685 ;
        RECT 0.900 3.455 1.420 3.635 ;
        RECT 1.090 2.975 1.420 3.455 ;
        RECT 1.610 2.975 1.940 3.805 ;
        RECT 0.000 2.635 0.920 2.805 ;
        RECT 0.095 1.495 0.425 2.635 ;
        RECT 1.090 2.465 1.295 2.975 ;
        RECT 2.135 2.805 2.465 3.975 ;
        RECT 2.660 3.935 3.360 3.975 ;
        RECT 2.660 3.805 3.140 3.935 ;
        RECT 2.660 2.975 2.990 3.805 ;
        RECT 3.530 3.685 3.700 4.435 ;
        RECT 5.040 4.435 5.430 4.605 ;
        RECT 5.600 4.685 6.040 4.855 ;
        RECT 6.275 4.780 6.605 5.355 ;
        RECT 6.840 4.855 7.090 5.110 ;
        RECT 6.840 4.685 7.280 4.855 ;
        RECT 3.305 3.635 3.700 3.685 ;
        RECT 3.180 3.455 3.700 3.635 ;
        RECT 3.180 2.975 3.510 3.455 ;
        RECT 1.465 2.635 3.135 2.805 ;
        RECT 1.090 1.985 1.420 2.465 ;
        RECT 0.900 1.805 1.420 1.985 ;
        RECT 0.900 1.755 1.295 1.805 ;
        RECT 0.900 1.005 1.070 1.755 ;
        RECT 1.610 1.635 1.940 2.465 ;
        RECT 1.460 1.505 1.940 1.635 ;
        RECT 1.240 1.465 1.940 1.505 ;
        RECT 2.135 1.465 2.465 2.635 ;
        RECT 3.305 2.465 3.510 2.975 ;
        RECT 4.175 2.805 4.565 3.945 ;
        RECT 5.040 3.685 5.210 4.435 ;
        RECT 5.600 4.265 5.770 4.685 ;
        RECT 5.380 3.975 5.770 4.265 ;
        RECT 7.110 4.265 7.280 4.685 ;
        RECT 7.450 4.605 7.695 5.110 ;
        RECT 7.450 4.435 7.840 4.605 ;
        RECT 8.350 4.555 8.670 5.355 ;
        RECT 9.325 4.605 9.570 5.110 ;
        RECT 9.930 4.855 10.180 5.110 ;
        RECT 7.110 3.975 7.500 4.265 ;
        RECT 5.380 3.935 6.080 3.975 ;
        RECT 5.600 3.805 6.080 3.935 ;
        RECT 5.040 3.635 5.435 3.685 ;
        RECT 5.040 3.455 5.560 3.635 ;
        RECT 5.230 2.975 5.560 3.455 ;
        RECT 5.750 2.975 6.080 3.805 ;
        RECT 3.680 2.635 5.060 2.805 ;
        RECT 2.660 1.635 2.990 2.465 ;
        RECT 3.180 1.985 3.510 2.465 ;
        RECT 3.180 1.805 3.700 1.985 ;
        RECT 3.305 1.755 3.700 1.805 ;
        RECT 2.660 1.505 3.140 1.635 ;
        RECT 2.660 1.465 3.360 1.505 ;
        RECT 1.240 1.175 1.630 1.465 ;
        RECT 0.130 0.085 0.390 0.885 ;
        RECT 0.900 0.835 1.290 1.005 ;
        RECT 1.045 0.330 1.290 0.835 ;
        RECT 1.460 0.755 1.630 1.175 ;
        RECT 2.970 1.175 3.360 1.465 ;
        RECT 2.970 0.755 3.140 1.175 ;
        RECT 3.530 1.005 3.700 1.755 ;
        RECT 4.175 1.495 4.565 2.635 ;
        RECT 5.230 2.465 5.435 2.975 ;
        RECT 6.275 2.805 6.605 3.975 ;
        RECT 6.800 3.935 7.500 3.975 ;
        RECT 6.800 3.805 7.280 3.935 ;
        RECT 6.800 2.975 7.130 3.805 ;
        RECT 7.670 3.685 7.840 4.435 ;
        RECT 9.180 4.435 9.570 4.605 ;
        RECT 9.740 4.685 10.180 4.855 ;
        RECT 10.415 4.780 10.745 5.355 ;
        RECT 10.980 4.855 11.230 5.110 ;
        RECT 10.980 4.685 11.420 4.855 ;
        RECT 7.445 3.635 7.840 3.685 ;
        RECT 7.320 3.455 7.840 3.635 ;
        RECT 7.320 2.975 7.650 3.455 ;
        RECT 5.605 2.635 7.275 2.805 ;
        RECT 5.230 1.985 5.560 2.465 ;
        RECT 5.040 1.805 5.560 1.985 ;
        RECT 5.040 1.755 5.435 1.805 ;
        RECT 1.460 0.585 1.900 0.755 ;
        RECT 1.650 0.330 1.900 0.585 ;
        RECT 2.135 0.085 2.465 0.660 ;
        RECT 2.700 0.585 3.140 0.755 ;
        RECT 3.310 0.835 3.700 1.005 ;
        RECT 5.040 1.005 5.210 1.755 ;
        RECT 5.750 1.635 6.080 2.465 ;
        RECT 5.600 1.505 6.080 1.635 ;
        RECT 5.380 1.465 6.080 1.505 ;
        RECT 6.275 1.465 6.605 2.635 ;
        RECT 7.445 2.465 7.650 2.975 ;
        RECT 8.315 2.805 8.705 3.945 ;
        RECT 9.180 3.685 9.350 4.435 ;
        RECT 9.740 4.265 9.910 4.685 ;
        RECT 9.520 3.975 9.910 4.265 ;
        RECT 11.250 4.265 11.420 4.685 ;
        RECT 11.590 4.605 11.835 5.110 ;
        RECT 11.590 4.435 11.980 4.605 ;
        RECT 12.490 4.555 12.810 5.355 ;
        RECT 13.465 4.605 13.710 5.110 ;
        RECT 14.070 4.855 14.320 5.110 ;
        RECT 11.250 3.975 11.640 4.265 ;
        RECT 9.520 3.935 10.220 3.975 ;
        RECT 9.740 3.805 10.220 3.935 ;
        RECT 9.180 3.635 9.575 3.685 ;
        RECT 9.180 3.455 9.700 3.635 ;
        RECT 9.370 2.975 9.700 3.455 ;
        RECT 9.890 2.975 10.220 3.805 ;
        RECT 7.820 2.635 9.200 2.805 ;
        RECT 6.800 1.635 7.130 2.465 ;
        RECT 7.320 1.985 7.650 2.465 ;
        RECT 7.320 1.805 7.840 1.985 ;
        RECT 7.445 1.755 7.840 1.805 ;
        RECT 6.800 1.505 7.280 1.635 ;
        RECT 6.800 1.465 7.500 1.505 ;
        RECT 5.380 1.175 5.770 1.465 ;
        RECT 2.700 0.330 2.950 0.585 ;
        RECT 3.310 0.330 3.555 0.835 ;
        RECT 4.210 0.085 4.530 0.885 ;
        RECT 5.040 0.835 5.430 1.005 ;
        RECT 5.185 0.330 5.430 0.835 ;
        RECT 5.600 0.755 5.770 1.175 ;
        RECT 7.110 1.175 7.500 1.465 ;
        RECT 7.110 0.755 7.280 1.175 ;
        RECT 7.670 1.005 7.840 1.755 ;
        RECT 8.315 1.495 8.705 2.635 ;
        RECT 9.370 2.465 9.575 2.975 ;
        RECT 10.415 2.805 10.745 3.975 ;
        RECT 10.940 3.935 11.640 3.975 ;
        RECT 10.940 3.805 11.420 3.935 ;
        RECT 10.940 2.975 11.270 3.805 ;
        RECT 11.810 3.685 11.980 4.435 ;
        RECT 13.320 4.435 13.710 4.605 ;
        RECT 13.880 4.685 14.320 4.855 ;
        RECT 14.555 4.780 14.885 5.355 ;
        RECT 15.120 4.855 15.370 5.110 ;
        RECT 15.120 4.685 15.560 4.855 ;
        RECT 11.585 3.635 11.980 3.685 ;
        RECT 11.460 3.455 11.980 3.635 ;
        RECT 11.460 2.975 11.790 3.455 ;
        RECT 9.745 2.635 11.415 2.805 ;
        RECT 9.370 1.985 9.700 2.465 ;
        RECT 9.180 1.805 9.700 1.985 ;
        RECT 9.180 1.755 9.575 1.805 ;
        RECT 5.600 0.585 6.040 0.755 ;
        RECT 5.790 0.330 6.040 0.585 ;
        RECT 6.275 0.085 6.605 0.660 ;
        RECT 6.840 0.585 7.280 0.755 ;
        RECT 7.450 0.835 7.840 1.005 ;
        RECT 9.180 1.005 9.350 1.755 ;
        RECT 9.890 1.635 10.220 2.465 ;
        RECT 9.740 1.505 10.220 1.635 ;
        RECT 9.520 1.465 10.220 1.505 ;
        RECT 10.415 1.465 10.745 2.635 ;
        RECT 11.585 2.465 11.790 2.975 ;
        RECT 12.455 2.805 12.845 3.945 ;
        RECT 13.320 3.685 13.490 4.435 ;
        RECT 13.880 4.265 14.050 4.685 ;
        RECT 13.660 3.975 14.050 4.265 ;
        RECT 15.390 4.265 15.560 4.685 ;
        RECT 15.730 4.605 15.975 5.110 ;
        RECT 15.730 4.435 16.120 4.605 ;
        RECT 16.630 4.555 16.890 5.355 ;
        RECT 15.390 3.975 15.780 4.265 ;
        RECT 13.660 3.935 14.360 3.975 ;
        RECT 13.880 3.805 14.360 3.935 ;
        RECT 13.320 3.635 13.715 3.685 ;
        RECT 13.320 3.455 13.840 3.635 ;
        RECT 13.510 2.975 13.840 3.455 ;
        RECT 14.030 2.975 14.360 3.805 ;
        RECT 11.960 2.635 13.340 2.805 ;
        RECT 10.940 1.635 11.270 2.465 ;
        RECT 11.460 1.985 11.790 2.465 ;
        RECT 11.460 1.805 11.980 1.985 ;
        RECT 11.585 1.755 11.980 1.805 ;
        RECT 10.940 1.505 11.420 1.635 ;
        RECT 10.940 1.465 11.640 1.505 ;
        RECT 9.520 1.175 9.910 1.465 ;
        RECT 6.840 0.330 7.090 0.585 ;
        RECT 7.450 0.330 7.695 0.835 ;
        RECT 8.350 0.085 8.670 0.885 ;
        RECT 9.180 0.835 9.570 1.005 ;
        RECT 9.325 0.330 9.570 0.835 ;
        RECT 9.740 0.755 9.910 1.175 ;
        RECT 11.250 1.175 11.640 1.465 ;
        RECT 11.250 0.755 11.420 1.175 ;
        RECT 11.810 1.005 11.980 1.755 ;
        RECT 12.455 1.495 12.845 2.635 ;
        RECT 13.510 2.465 13.715 2.975 ;
        RECT 14.555 2.805 14.885 3.975 ;
        RECT 15.080 3.935 15.780 3.975 ;
        RECT 15.080 3.805 15.560 3.935 ;
        RECT 15.080 2.975 15.410 3.805 ;
        RECT 15.950 3.685 16.120 4.435 ;
        RECT 15.725 3.635 16.120 3.685 ;
        RECT 15.600 3.455 16.120 3.635 ;
        RECT 15.600 2.975 15.930 3.455 ;
        RECT 13.885 2.635 15.555 2.805 ;
        RECT 13.510 1.985 13.840 2.465 ;
        RECT 13.320 1.805 13.840 1.985 ;
        RECT 13.320 1.755 13.715 1.805 ;
        RECT 9.740 0.585 10.180 0.755 ;
        RECT 9.930 0.330 10.180 0.585 ;
        RECT 10.415 0.085 10.745 0.660 ;
        RECT 10.980 0.585 11.420 0.755 ;
        RECT 11.590 0.835 11.980 1.005 ;
        RECT 13.320 1.005 13.490 1.755 ;
        RECT 14.030 1.635 14.360 2.465 ;
        RECT 13.880 1.505 14.360 1.635 ;
        RECT 13.660 1.465 14.360 1.505 ;
        RECT 14.555 1.465 14.885 2.635 ;
        RECT 15.725 2.465 15.930 2.975 ;
        RECT 16.595 2.805 16.925 3.945 ;
        RECT 16.100 2.635 17.020 2.805 ;
        RECT 15.080 1.635 15.410 2.465 ;
        RECT 15.600 1.985 15.930 2.465 ;
        RECT 15.600 1.805 16.120 1.985 ;
        RECT 15.725 1.755 16.120 1.805 ;
        RECT 15.080 1.505 15.560 1.635 ;
        RECT 15.080 1.465 15.780 1.505 ;
        RECT 13.660 1.175 14.050 1.465 ;
        RECT 10.980 0.330 11.230 0.585 ;
        RECT 11.590 0.330 11.835 0.835 ;
        RECT 12.490 0.085 12.810 0.885 ;
        RECT 13.320 0.835 13.710 1.005 ;
        RECT 13.465 0.330 13.710 0.835 ;
        RECT 13.880 0.755 14.050 1.175 ;
        RECT 15.390 1.175 15.780 1.465 ;
        RECT 15.390 0.755 15.560 1.175 ;
        RECT 15.950 1.005 16.120 1.755 ;
        RECT 16.595 1.495 16.925 2.635 ;
        RECT 13.880 0.585 14.320 0.755 ;
        RECT 14.070 0.330 14.320 0.585 ;
        RECT 14.555 0.085 14.885 0.660 ;
        RECT 15.120 0.585 15.560 0.755 ;
        RECT 15.730 0.835 16.120 1.005 ;
        RECT 15.120 0.330 15.370 0.585 ;
        RECT 15.730 0.330 15.975 0.835 ;
        RECT 16.630 0.085 16.890 0.885 ;
        RECT 0.000 -0.085 17.020 0.085 ;
      LAYER mcon ;
        RECT 0.145 5.355 0.315 5.525 ;
        RECT 0.605 5.355 0.775 5.525 ;
        RECT 1.065 5.355 1.235 5.525 ;
        RECT 1.525 5.355 1.695 5.525 ;
        RECT 1.985 5.355 2.155 5.525 ;
        RECT 2.445 5.355 2.615 5.525 ;
        RECT 2.905 5.355 3.075 5.525 ;
        RECT 3.365 5.355 3.535 5.525 ;
        RECT 3.825 5.355 3.995 5.525 ;
        RECT 4.285 5.355 4.455 5.525 ;
        RECT 4.745 5.355 4.915 5.525 ;
        RECT 5.205 5.355 5.375 5.525 ;
        RECT 5.665 5.355 5.835 5.525 ;
        RECT 6.125 5.355 6.295 5.525 ;
        RECT 6.585 5.355 6.755 5.525 ;
        RECT 7.045 5.355 7.215 5.525 ;
        RECT 7.505 5.355 7.675 5.525 ;
        RECT 7.965 5.355 8.135 5.525 ;
        RECT 8.425 5.355 8.595 5.525 ;
        RECT 8.885 5.355 9.055 5.525 ;
        RECT 9.345 5.355 9.515 5.525 ;
        RECT 9.805 5.355 9.975 5.525 ;
        RECT 10.265 5.355 10.435 5.525 ;
        RECT 10.725 5.355 10.895 5.525 ;
        RECT 11.185 5.355 11.355 5.525 ;
        RECT 11.645 5.355 11.815 5.525 ;
        RECT 12.105 5.355 12.275 5.525 ;
        RECT 12.565 5.355 12.735 5.525 ;
        RECT 13.025 5.355 13.195 5.525 ;
        RECT 13.485 5.355 13.655 5.525 ;
        RECT 13.945 5.355 14.115 5.525 ;
        RECT 14.405 5.355 14.575 5.525 ;
        RECT 14.865 5.355 15.035 5.525 ;
        RECT 15.325 5.355 15.495 5.525 ;
        RECT 15.785 5.355 15.955 5.525 ;
        RECT 16.245 5.355 16.415 5.525 ;
        RECT 16.705 5.355 16.875 5.525 ;
        RECT 1.065 3.485 1.235 3.655 ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 3.365 3.485 3.535 3.655 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 1.065 1.785 1.235 1.955 ;
        RECT 5.205 3.485 5.375 3.655 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 3.365 1.785 3.535 1.955 ;
        RECT 7.505 3.485 7.675 3.655 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 5.205 1.785 5.375 1.955 ;
        RECT 9.345 3.485 9.515 3.655 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 7.505 1.785 7.675 1.955 ;
        RECT 11.645 3.485 11.815 3.655 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 9.345 1.785 9.515 1.955 ;
        RECT 13.485 3.485 13.655 3.655 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 11.645 1.785 11.815 1.955 ;
        RECT 15.785 3.485 15.955 3.655 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 14.405 2.635 14.575 2.805 ;
        RECT 14.865 2.635 15.035 2.805 ;
        RECT 15.325 2.635 15.495 2.805 ;
        RECT 13.485 1.785 13.655 1.955 ;
        RECT 16.245 2.635 16.415 2.805 ;
        RECT 16.705 2.635 16.875 2.805 ;
        RECT 15.785 1.785 15.955 1.955 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
        RECT 14.405 -0.085 14.575 0.085 ;
        RECT 14.865 -0.085 15.035 0.085 ;
        RECT 15.325 -0.085 15.495 0.085 ;
        RECT 15.785 -0.085 15.955 0.085 ;
        RECT 16.245 -0.085 16.415 0.085 ;
        RECT 16.705 -0.085 16.875 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__muxb16to1_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__muxb16to1_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__muxb16to1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.760 BY 5.440 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 24.845 4.115 25.665 4.385 ;
    END
  END D[15]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 19.415 4.115 20.235 4.385 ;
    END
  END D[14]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 18.405 4.115 19.225 4.385 ;
    END
  END D[13]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 12.975 4.115 13.795 4.385 ;
    END
  END D[12]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 11.965 4.115 12.785 4.385 ;
    END
  END D[11]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 6.535 4.115 7.355 4.385 ;
    END
  END D[10]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 5.525 4.115 6.345 4.385 ;
    END
  END D[9]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.095 4.115 0.915 4.385 ;
    END
  END D[8]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 24.845 1.055 25.665 1.325 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 19.415 1.055 20.235 1.325 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 18.405 1.055 19.225 1.325 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 12.975 1.055 13.795 1.325 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 11.965 1.055 12.785 1.325 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 6.535 1.055 7.355 1.325 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 5.525 1.055 6.345 1.325 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.055 0.915 1.325 ;
    END
  END D[0]
  PIN S[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 22.635 4.145 22.970 4.415 ;
    END
  END S[15]
  PIN S[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 22.110 4.145 22.445 4.415 ;
    END
  END S[14]
  PIN S[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 16.195 4.145 16.530 4.415 ;
    END
  END S[13]
  PIN S[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 15.670 4.145 16.005 4.415 ;
    END
  END S[12]
  PIN S[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 9.755 4.145 10.090 4.415 ;
    END
  END S[11]
  PIN S[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 9.230 4.145 9.565 4.415 ;
    END
  END S[10]
  PIN S[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 3.315 4.145 3.650 4.415 ;
    END
  END S[9]
  PIN S[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 2.790 4.145 3.125 4.415 ;
    END
  END S[8]
  PIN S[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 22.635 1.025 22.970 1.295 ;
    END
  END S[7]
  PIN S[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 22.110 1.025 22.445 1.295 ;
    END
  END S[6]
  PIN S[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 16.195 1.025 16.530 1.295 ;
    END
  END S[5]
  PIN S[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 15.670 1.025 16.005 1.295 ;
    END
  END S[4]
  PIN S[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 9.755 1.025 10.090 1.295 ;
    END
  END S[3]
  PIN S[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 9.230 1.025 9.565 1.295 ;
    END
  END S[2]
  PIN S[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 3.315 1.025 3.650 1.295 ;
    END
  END S[1]
  PIN S[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 2.790 1.025 3.125 1.295 ;
    END
  END S[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 25.760 0.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 5.200 25.760 5.680 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.995 1.440 1.015 ;
        RECT 5.000 0.995 7.880 1.015 ;
        RECT 11.440 0.995 14.320 1.015 ;
        RECT 17.880 0.995 20.760 1.015 ;
        RECT 24.320 0.995 25.755 1.015 ;
        RECT 0.005 0.885 2.345 0.995 ;
        RECT 4.095 0.885 8.785 0.995 ;
        RECT 10.535 0.885 15.225 0.995 ;
        RECT 16.975 0.885 21.665 0.995 ;
        RECT 23.415 0.885 25.755 0.995 ;
        RECT 0.005 0.215 25.755 0.885 ;
        RECT 0.005 0.105 1.440 0.215 ;
        RECT 2.545 0.105 3.895 0.215 ;
        RECT 5.000 0.105 7.880 0.215 ;
        RECT 8.985 0.105 10.335 0.215 ;
        RECT 11.440 0.105 14.320 0.215 ;
        RECT 15.425 0.105 16.775 0.215 ;
        RECT 17.880 0.105 20.760 0.215 ;
        RECT 21.865 0.105 23.215 0.215 ;
        RECT 24.320 0.105 25.755 0.215 ;
        RECT 0.145 -0.085 0.315 0.105 ;
        RECT 6.125 -0.085 6.755 0.105 ;
        RECT 12.565 -0.085 13.195 0.105 ;
        RECT 19.005 -0.085 19.635 0.105 ;
        RECT 25.445 -0.085 25.615 0.105 ;
    END
    PORT
      LAYER pwell ;
        RECT 0.145 5.335 0.315 5.525 ;
        RECT 6.125 5.335 6.755 5.525 ;
        RECT 12.565 5.335 13.195 5.525 ;
        RECT 19.005 5.335 19.635 5.525 ;
        RECT 25.445 5.335 25.615 5.525 ;
        RECT 0.005 5.225 1.440 5.335 ;
        RECT 2.545 5.225 3.895 5.335 ;
        RECT 5.000 5.225 7.880 5.335 ;
        RECT 8.985 5.225 10.335 5.335 ;
        RECT 11.440 5.225 14.320 5.335 ;
        RECT 15.425 5.225 16.775 5.335 ;
        RECT 17.880 5.225 20.760 5.335 ;
        RECT 21.865 5.225 23.215 5.335 ;
        RECT 24.320 5.225 25.755 5.335 ;
        RECT 0.005 4.555 25.755 5.225 ;
        RECT 0.005 4.445 2.345 4.555 ;
        RECT 4.095 4.445 8.785 4.555 ;
        RECT 10.535 4.445 15.225 4.555 ;
        RECT 16.975 4.445 21.665 4.555 ;
        RECT 23.415 4.445 25.755 4.555 ;
        RECT 0.005 4.425 1.440 4.445 ;
        RECT 5.000 4.425 7.880 4.445 ;
        RECT 11.440 4.425 14.320 4.445 ;
        RECT 17.880 4.425 20.760 4.445 ;
        RECT 24.320 4.425 25.755 4.445 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 25.950 4.135 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 25.760 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.051200 ;
    PORT
      LAYER met1 ;
        RECT 1.465 3.640 1.755 3.685 ;
        RECT 4.685 3.640 4.975 3.685 ;
        RECT 7.905 3.640 8.195 3.685 ;
        RECT 11.125 3.640 11.415 3.685 ;
        RECT 14.345 3.640 14.635 3.685 ;
        RECT 17.565 3.640 17.855 3.685 ;
        RECT 20.785 3.640 21.075 3.685 ;
        RECT 24.005 3.640 24.295 3.685 ;
        RECT 1.465 3.500 24.295 3.640 ;
        RECT 1.465 3.455 1.755 3.500 ;
        RECT 4.685 3.455 4.975 3.500 ;
        RECT 7.905 3.455 8.195 3.500 ;
        RECT 11.125 3.455 11.415 3.500 ;
        RECT 14.345 3.455 14.635 3.500 ;
        RECT 17.565 3.455 17.855 3.500 ;
        RECT 20.785 3.455 21.075 3.500 ;
        RECT 24.005 3.455 24.295 3.500 ;
        RECT 1.465 1.940 1.755 1.985 ;
        RECT 4.685 1.940 4.975 1.985 ;
        RECT 7.905 1.940 8.195 1.985 ;
        RECT 11.125 1.940 11.415 1.985 ;
        RECT 14.345 1.940 14.635 1.985 ;
        RECT 17.565 1.940 17.855 1.985 ;
        RECT 20.785 1.940 21.075 1.985 ;
        RECT 24.005 1.940 24.295 1.985 ;
        RECT 1.465 1.800 24.295 1.940 ;
        RECT 1.465 1.755 1.755 1.800 ;
        RECT 4.685 1.755 4.975 1.800 ;
        RECT 7.905 1.755 8.195 1.800 ;
        RECT 11.125 1.755 11.415 1.800 ;
        RECT 14.345 1.755 14.635 1.800 ;
        RECT 17.565 1.755 17.855 1.800 ;
        RECT 20.785 1.755 21.075 1.800 ;
        RECT 24.005 1.755 24.295 1.800 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 5.355 25.760 5.525 ;
        RECT 0.145 4.725 0.475 5.185 ;
        RECT 0.645 4.895 0.860 5.355 ;
        RECT 1.030 5.015 2.175 5.185 ;
        RECT 1.030 4.725 1.335 5.015 ;
        RECT 0.145 4.555 1.335 4.725 ;
        RECT 1.505 4.555 1.835 4.845 ;
        RECT 2.005 4.670 2.175 5.015 ;
        RECT 2.675 4.855 2.925 5.110 ;
        RECT 2.345 4.685 2.925 4.855 ;
        RECT 3.095 4.780 3.345 5.355 ;
        RECT 3.515 4.855 3.765 5.110 ;
        RECT 4.265 5.015 5.410 5.185 ;
        RECT 3.515 4.685 4.095 4.855 ;
        RECT 1.030 4.515 1.335 4.555 ;
        RECT 0.095 3.775 1.285 3.945 ;
        RECT 0.095 3.230 0.395 3.775 ;
        RECT 0.565 3.335 0.895 3.605 ;
        RECT 0.095 2.975 0.425 3.230 ;
        RECT 0.595 2.805 0.895 3.335 ;
        RECT 1.115 3.145 1.285 3.775 ;
        RECT 1.585 3.685 1.755 4.555 ;
        RECT 2.345 4.235 2.515 4.685 ;
        RECT 2.100 4.135 2.515 4.235 ;
        RECT 3.925 4.235 4.095 4.685 ;
        RECT 4.265 4.670 4.435 5.015 ;
        RECT 4.605 4.555 4.935 4.845 ;
        RECT 5.105 4.725 5.410 5.015 ;
        RECT 5.580 4.895 5.795 5.355 ;
        RECT 5.965 4.725 6.295 5.185 ;
        RECT 5.105 4.555 6.295 4.725 ;
        RECT 6.585 4.725 6.915 5.185 ;
        RECT 7.085 4.895 7.300 5.355 ;
        RECT 7.470 5.015 8.615 5.185 ;
        RECT 7.470 4.725 7.775 5.015 ;
        RECT 6.585 4.555 7.775 4.725 ;
        RECT 7.945 4.555 8.275 4.845 ;
        RECT 8.445 4.670 8.615 5.015 ;
        RECT 9.115 4.855 9.365 5.110 ;
        RECT 8.785 4.685 9.365 4.855 ;
        RECT 9.535 4.780 9.785 5.355 ;
        RECT 9.955 4.855 10.205 5.110 ;
        RECT 10.705 5.015 11.850 5.185 ;
        RECT 9.955 4.685 10.535 4.855 ;
        RECT 3.925 4.135 4.340 4.235 ;
        RECT 2.100 3.975 2.620 4.135 ;
        RECT 3.820 3.975 4.340 4.135 ;
        RECT 2.100 3.965 2.880 3.975 ;
        RECT 2.450 3.805 2.880 3.965 ;
        RECT 1.465 3.315 1.895 3.685 ;
        RECT 1.115 2.975 1.415 3.145 ;
        RECT 0.000 2.635 1.415 2.805 ;
        RECT 0.095 2.210 0.425 2.465 ;
        RECT 0.095 1.665 0.395 2.210 ;
        RECT 0.595 2.105 0.895 2.635 ;
        RECT 0.565 1.835 0.895 2.105 ;
        RECT 1.115 2.295 1.415 2.465 ;
        RECT 1.115 1.665 1.285 2.295 ;
        RECT 1.585 2.125 1.755 3.315 ;
        RECT 2.110 3.145 2.280 3.795 ;
        RECT 1.925 2.975 2.280 3.145 ;
        RECT 2.550 2.975 2.880 3.805 ;
        RECT 3.055 2.805 3.385 3.975 ;
        RECT 3.560 3.965 4.340 3.975 ;
        RECT 3.560 3.805 3.990 3.965 ;
        RECT 3.560 2.975 3.890 3.805 ;
        RECT 4.160 3.145 4.330 3.795 ;
        RECT 4.685 3.685 4.855 4.555 ;
        RECT 5.105 4.515 5.410 4.555 ;
        RECT 7.470 4.515 7.775 4.555 ;
        RECT 5.155 3.775 6.345 3.945 ;
        RECT 4.545 3.315 4.975 3.685 ;
        RECT 4.160 2.975 4.515 3.145 ;
        RECT 1.925 2.635 4.515 2.805 ;
        RECT 1.925 2.295 2.280 2.465 ;
        RECT 1.465 1.755 1.895 2.125 ;
        RECT 0.095 1.495 1.285 1.665 ;
        RECT 1.030 0.885 1.335 0.925 ;
        RECT 1.585 0.885 1.755 1.755 ;
        RECT 2.110 1.645 2.280 2.295 ;
        RECT 2.550 1.635 2.880 2.465 ;
        RECT 2.450 1.475 2.880 1.635 ;
        RECT 2.100 1.465 2.880 1.475 ;
        RECT 3.055 1.465 3.385 2.635 ;
        RECT 3.560 1.635 3.890 2.465 ;
        RECT 4.160 2.295 4.515 2.465 ;
        RECT 4.160 1.645 4.330 2.295 ;
        RECT 4.685 2.125 4.855 3.315 ;
        RECT 5.155 3.145 5.325 3.775 ;
        RECT 5.025 2.975 5.325 3.145 ;
        RECT 5.545 3.335 5.875 3.605 ;
        RECT 5.545 2.805 5.845 3.335 ;
        RECT 6.045 3.230 6.345 3.775 ;
        RECT 6.015 2.975 6.345 3.230 ;
        RECT 6.535 3.775 7.725 3.945 ;
        RECT 6.535 3.230 6.835 3.775 ;
        RECT 7.005 3.335 7.335 3.605 ;
        RECT 6.535 2.975 6.865 3.230 ;
        RECT 7.035 2.805 7.335 3.335 ;
        RECT 7.555 3.145 7.725 3.775 ;
        RECT 8.025 3.685 8.195 4.555 ;
        RECT 8.785 4.235 8.955 4.685 ;
        RECT 8.540 4.135 8.955 4.235 ;
        RECT 10.365 4.235 10.535 4.685 ;
        RECT 10.705 4.670 10.875 5.015 ;
        RECT 11.045 4.555 11.375 4.845 ;
        RECT 11.545 4.725 11.850 5.015 ;
        RECT 12.020 4.895 12.235 5.355 ;
        RECT 12.405 4.725 12.735 5.185 ;
        RECT 11.545 4.555 12.735 4.725 ;
        RECT 13.025 4.725 13.355 5.185 ;
        RECT 13.525 4.895 13.740 5.355 ;
        RECT 13.910 5.015 15.055 5.185 ;
        RECT 13.910 4.725 14.215 5.015 ;
        RECT 13.025 4.555 14.215 4.725 ;
        RECT 14.385 4.555 14.715 4.845 ;
        RECT 14.885 4.670 15.055 5.015 ;
        RECT 15.555 4.855 15.805 5.110 ;
        RECT 15.225 4.685 15.805 4.855 ;
        RECT 15.975 4.780 16.225 5.355 ;
        RECT 16.395 4.855 16.645 5.110 ;
        RECT 17.145 5.015 18.290 5.185 ;
        RECT 16.395 4.685 16.975 4.855 ;
        RECT 10.365 4.135 10.780 4.235 ;
        RECT 8.540 3.975 9.060 4.135 ;
        RECT 10.260 3.975 10.780 4.135 ;
        RECT 8.540 3.965 9.320 3.975 ;
        RECT 8.890 3.805 9.320 3.965 ;
        RECT 7.905 3.315 8.335 3.685 ;
        RECT 7.555 2.975 7.855 3.145 ;
        RECT 5.025 2.635 7.855 2.805 ;
        RECT 5.025 2.295 5.325 2.465 ;
        RECT 4.545 1.755 4.975 2.125 ;
        RECT 3.560 1.475 3.990 1.635 ;
        RECT 3.560 1.465 4.340 1.475 ;
        RECT 2.100 1.305 2.620 1.465 ;
        RECT 3.820 1.305 4.340 1.465 ;
        RECT 2.100 1.205 2.515 1.305 ;
        RECT 0.145 0.715 1.335 0.885 ;
        RECT 0.145 0.255 0.475 0.715 ;
        RECT 0.645 0.085 0.860 0.545 ;
        RECT 1.030 0.425 1.335 0.715 ;
        RECT 1.505 0.595 1.835 0.885 ;
        RECT 2.005 0.425 2.175 0.770 ;
        RECT 2.345 0.755 2.515 1.205 ;
        RECT 3.925 1.205 4.340 1.305 ;
        RECT 3.925 0.755 4.095 1.205 ;
        RECT 4.685 0.885 4.855 1.755 ;
        RECT 5.155 1.665 5.325 2.295 ;
        RECT 5.545 2.105 5.845 2.635 ;
        RECT 6.015 2.210 6.345 2.465 ;
        RECT 5.545 1.835 5.875 2.105 ;
        RECT 6.045 1.665 6.345 2.210 ;
        RECT 5.155 1.495 6.345 1.665 ;
        RECT 6.535 2.210 6.865 2.465 ;
        RECT 6.535 1.665 6.835 2.210 ;
        RECT 7.035 2.105 7.335 2.635 ;
        RECT 7.005 1.835 7.335 2.105 ;
        RECT 7.555 2.295 7.855 2.465 ;
        RECT 7.555 1.665 7.725 2.295 ;
        RECT 8.025 2.125 8.195 3.315 ;
        RECT 8.550 3.145 8.720 3.795 ;
        RECT 8.365 2.975 8.720 3.145 ;
        RECT 8.990 2.975 9.320 3.805 ;
        RECT 9.495 2.805 9.825 3.975 ;
        RECT 10.000 3.965 10.780 3.975 ;
        RECT 10.000 3.805 10.430 3.965 ;
        RECT 10.000 2.975 10.330 3.805 ;
        RECT 10.600 3.145 10.770 3.795 ;
        RECT 11.125 3.685 11.295 4.555 ;
        RECT 11.545 4.515 11.850 4.555 ;
        RECT 13.910 4.515 14.215 4.555 ;
        RECT 11.595 3.775 12.785 3.945 ;
        RECT 10.985 3.315 11.415 3.685 ;
        RECT 10.600 2.975 10.955 3.145 ;
        RECT 8.365 2.635 10.955 2.805 ;
        RECT 8.365 2.295 8.720 2.465 ;
        RECT 7.905 1.755 8.335 2.125 ;
        RECT 6.535 1.495 7.725 1.665 ;
        RECT 5.105 0.885 5.410 0.925 ;
        RECT 7.470 0.885 7.775 0.925 ;
        RECT 8.025 0.885 8.195 1.755 ;
        RECT 8.550 1.645 8.720 2.295 ;
        RECT 8.990 1.635 9.320 2.465 ;
        RECT 8.890 1.475 9.320 1.635 ;
        RECT 8.540 1.465 9.320 1.475 ;
        RECT 9.495 1.465 9.825 2.635 ;
        RECT 10.000 1.635 10.330 2.465 ;
        RECT 10.600 2.295 10.955 2.465 ;
        RECT 10.600 1.645 10.770 2.295 ;
        RECT 11.125 2.125 11.295 3.315 ;
        RECT 11.595 3.145 11.765 3.775 ;
        RECT 11.465 2.975 11.765 3.145 ;
        RECT 11.985 3.335 12.315 3.605 ;
        RECT 11.985 2.805 12.285 3.335 ;
        RECT 12.485 3.230 12.785 3.775 ;
        RECT 12.455 2.975 12.785 3.230 ;
        RECT 12.975 3.775 14.165 3.945 ;
        RECT 12.975 3.230 13.275 3.775 ;
        RECT 13.445 3.335 13.775 3.605 ;
        RECT 12.975 2.975 13.305 3.230 ;
        RECT 13.475 2.805 13.775 3.335 ;
        RECT 13.995 3.145 14.165 3.775 ;
        RECT 14.465 3.685 14.635 4.555 ;
        RECT 15.225 4.235 15.395 4.685 ;
        RECT 14.980 4.135 15.395 4.235 ;
        RECT 16.805 4.235 16.975 4.685 ;
        RECT 17.145 4.670 17.315 5.015 ;
        RECT 17.485 4.555 17.815 4.845 ;
        RECT 17.985 4.725 18.290 5.015 ;
        RECT 18.460 4.895 18.675 5.355 ;
        RECT 18.845 4.725 19.175 5.185 ;
        RECT 17.985 4.555 19.175 4.725 ;
        RECT 19.465 4.725 19.795 5.185 ;
        RECT 19.965 4.895 20.180 5.355 ;
        RECT 20.350 5.015 21.495 5.185 ;
        RECT 20.350 4.725 20.655 5.015 ;
        RECT 19.465 4.555 20.655 4.725 ;
        RECT 20.825 4.555 21.155 4.845 ;
        RECT 21.325 4.670 21.495 5.015 ;
        RECT 21.995 4.855 22.245 5.110 ;
        RECT 21.665 4.685 22.245 4.855 ;
        RECT 22.415 4.780 22.665 5.355 ;
        RECT 22.835 4.855 23.085 5.110 ;
        RECT 23.585 5.015 24.730 5.185 ;
        RECT 22.835 4.685 23.415 4.855 ;
        RECT 16.805 4.135 17.220 4.235 ;
        RECT 14.980 3.975 15.500 4.135 ;
        RECT 16.700 3.975 17.220 4.135 ;
        RECT 14.980 3.965 15.760 3.975 ;
        RECT 15.330 3.805 15.760 3.965 ;
        RECT 14.345 3.315 14.775 3.685 ;
        RECT 13.995 2.975 14.295 3.145 ;
        RECT 11.465 2.635 14.295 2.805 ;
        RECT 11.465 2.295 11.765 2.465 ;
        RECT 10.985 1.755 11.415 2.125 ;
        RECT 10.000 1.475 10.430 1.635 ;
        RECT 10.000 1.465 10.780 1.475 ;
        RECT 8.540 1.305 9.060 1.465 ;
        RECT 10.260 1.305 10.780 1.465 ;
        RECT 8.540 1.205 8.955 1.305 ;
        RECT 2.345 0.585 2.925 0.755 ;
        RECT 1.030 0.255 2.175 0.425 ;
        RECT 2.675 0.330 2.925 0.585 ;
        RECT 3.095 0.085 3.345 0.660 ;
        RECT 3.515 0.585 4.095 0.755 ;
        RECT 3.515 0.330 3.765 0.585 ;
        RECT 4.265 0.425 4.435 0.770 ;
        RECT 4.605 0.595 4.935 0.885 ;
        RECT 5.105 0.715 6.295 0.885 ;
        RECT 5.105 0.425 5.410 0.715 ;
        RECT 4.265 0.255 5.410 0.425 ;
        RECT 5.580 0.085 5.795 0.545 ;
        RECT 5.965 0.255 6.295 0.715 ;
        RECT 6.585 0.715 7.775 0.885 ;
        RECT 6.585 0.255 6.915 0.715 ;
        RECT 7.085 0.085 7.300 0.545 ;
        RECT 7.470 0.425 7.775 0.715 ;
        RECT 7.945 0.595 8.275 0.885 ;
        RECT 8.445 0.425 8.615 0.770 ;
        RECT 8.785 0.755 8.955 1.205 ;
        RECT 10.365 1.205 10.780 1.305 ;
        RECT 10.365 0.755 10.535 1.205 ;
        RECT 11.125 0.885 11.295 1.755 ;
        RECT 11.595 1.665 11.765 2.295 ;
        RECT 11.985 2.105 12.285 2.635 ;
        RECT 12.455 2.210 12.785 2.465 ;
        RECT 11.985 1.835 12.315 2.105 ;
        RECT 12.485 1.665 12.785 2.210 ;
        RECT 11.595 1.495 12.785 1.665 ;
        RECT 12.975 2.210 13.305 2.465 ;
        RECT 12.975 1.665 13.275 2.210 ;
        RECT 13.475 2.105 13.775 2.635 ;
        RECT 13.445 1.835 13.775 2.105 ;
        RECT 13.995 2.295 14.295 2.465 ;
        RECT 13.995 1.665 14.165 2.295 ;
        RECT 14.465 2.125 14.635 3.315 ;
        RECT 14.990 3.145 15.160 3.795 ;
        RECT 14.805 2.975 15.160 3.145 ;
        RECT 15.430 2.975 15.760 3.805 ;
        RECT 15.935 2.805 16.265 3.975 ;
        RECT 16.440 3.965 17.220 3.975 ;
        RECT 16.440 3.805 16.870 3.965 ;
        RECT 16.440 2.975 16.770 3.805 ;
        RECT 17.040 3.145 17.210 3.795 ;
        RECT 17.565 3.685 17.735 4.555 ;
        RECT 17.985 4.515 18.290 4.555 ;
        RECT 20.350 4.515 20.655 4.555 ;
        RECT 18.035 3.775 19.225 3.945 ;
        RECT 17.425 3.315 17.855 3.685 ;
        RECT 17.040 2.975 17.395 3.145 ;
        RECT 14.805 2.635 17.395 2.805 ;
        RECT 14.805 2.295 15.160 2.465 ;
        RECT 14.345 1.755 14.775 2.125 ;
        RECT 12.975 1.495 14.165 1.665 ;
        RECT 11.545 0.885 11.850 0.925 ;
        RECT 13.910 0.885 14.215 0.925 ;
        RECT 14.465 0.885 14.635 1.755 ;
        RECT 14.990 1.645 15.160 2.295 ;
        RECT 15.430 1.635 15.760 2.465 ;
        RECT 15.330 1.475 15.760 1.635 ;
        RECT 14.980 1.465 15.760 1.475 ;
        RECT 15.935 1.465 16.265 2.635 ;
        RECT 16.440 1.635 16.770 2.465 ;
        RECT 17.040 2.295 17.395 2.465 ;
        RECT 17.040 1.645 17.210 2.295 ;
        RECT 17.565 2.125 17.735 3.315 ;
        RECT 18.035 3.145 18.205 3.775 ;
        RECT 17.905 2.975 18.205 3.145 ;
        RECT 18.425 3.335 18.755 3.605 ;
        RECT 18.425 2.805 18.725 3.335 ;
        RECT 18.925 3.230 19.225 3.775 ;
        RECT 18.895 2.975 19.225 3.230 ;
        RECT 19.415 3.775 20.605 3.945 ;
        RECT 19.415 3.230 19.715 3.775 ;
        RECT 19.885 3.335 20.215 3.605 ;
        RECT 19.415 2.975 19.745 3.230 ;
        RECT 19.915 2.805 20.215 3.335 ;
        RECT 20.435 3.145 20.605 3.775 ;
        RECT 20.905 3.685 21.075 4.555 ;
        RECT 21.665 4.235 21.835 4.685 ;
        RECT 21.420 4.135 21.835 4.235 ;
        RECT 23.245 4.235 23.415 4.685 ;
        RECT 23.585 4.670 23.755 5.015 ;
        RECT 23.925 4.555 24.255 4.845 ;
        RECT 24.425 4.725 24.730 5.015 ;
        RECT 24.900 4.895 25.115 5.355 ;
        RECT 25.285 4.725 25.615 5.185 ;
        RECT 24.425 4.555 25.615 4.725 ;
        RECT 23.245 4.135 23.660 4.235 ;
        RECT 21.420 3.975 21.940 4.135 ;
        RECT 23.140 3.975 23.660 4.135 ;
        RECT 21.420 3.965 22.200 3.975 ;
        RECT 21.770 3.805 22.200 3.965 ;
        RECT 20.785 3.315 21.215 3.685 ;
        RECT 20.435 2.975 20.735 3.145 ;
        RECT 17.905 2.635 20.735 2.805 ;
        RECT 17.905 2.295 18.205 2.465 ;
        RECT 17.425 1.755 17.855 2.125 ;
        RECT 16.440 1.475 16.870 1.635 ;
        RECT 16.440 1.465 17.220 1.475 ;
        RECT 14.980 1.305 15.500 1.465 ;
        RECT 16.700 1.305 17.220 1.465 ;
        RECT 14.980 1.205 15.395 1.305 ;
        RECT 8.785 0.585 9.365 0.755 ;
        RECT 7.470 0.255 8.615 0.425 ;
        RECT 9.115 0.330 9.365 0.585 ;
        RECT 9.535 0.085 9.785 0.660 ;
        RECT 9.955 0.585 10.535 0.755 ;
        RECT 9.955 0.330 10.205 0.585 ;
        RECT 10.705 0.425 10.875 0.770 ;
        RECT 11.045 0.595 11.375 0.885 ;
        RECT 11.545 0.715 12.735 0.885 ;
        RECT 11.545 0.425 11.850 0.715 ;
        RECT 10.705 0.255 11.850 0.425 ;
        RECT 12.020 0.085 12.235 0.545 ;
        RECT 12.405 0.255 12.735 0.715 ;
        RECT 13.025 0.715 14.215 0.885 ;
        RECT 13.025 0.255 13.355 0.715 ;
        RECT 13.525 0.085 13.740 0.545 ;
        RECT 13.910 0.425 14.215 0.715 ;
        RECT 14.385 0.595 14.715 0.885 ;
        RECT 14.885 0.425 15.055 0.770 ;
        RECT 15.225 0.755 15.395 1.205 ;
        RECT 16.805 1.205 17.220 1.305 ;
        RECT 16.805 0.755 16.975 1.205 ;
        RECT 17.565 0.885 17.735 1.755 ;
        RECT 18.035 1.665 18.205 2.295 ;
        RECT 18.425 2.105 18.725 2.635 ;
        RECT 18.895 2.210 19.225 2.465 ;
        RECT 18.425 1.835 18.755 2.105 ;
        RECT 18.925 1.665 19.225 2.210 ;
        RECT 18.035 1.495 19.225 1.665 ;
        RECT 19.415 2.210 19.745 2.465 ;
        RECT 19.415 1.665 19.715 2.210 ;
        RECT 19.915 2.105 20.215 2.635 ;
        RECT 19.885 1.835 20.215 2.105 ;
        RECT 20.435 2.295 20.735 2.465 ;
        RECT 20.435 1.665 20.605 2.295 ;
        RECT 20.905 2.125 21.075 3.315 ;
        RECT 21.430 3.145 21.600 3.795 ;
        RECT 21.245 2.975 21.600 3.145 ;
        RECT 21.870 2.975 22.200 3.805 ;
        RECT 22.375 2.805 22.705 3.975 ;
        RECT 22.880 3.965 23.660 3.975 ;
        RECT 22.880 3.805 23.310 3.965 ;
        RECT 22.880 2.975 23.210 3.805 ;
        RECT 23.480 3.145 23.650 3.795 ;
        RECT 24.005 3.685 24.175 4.555 ;
        RECT 24.425 4.515 24.730 4.555 ;
        RECT 24.475 3.775 25.665 3.945 ;
        RECT 23.865 3.315 24.295 3.685 ;
        RECT 23.480 2.975 23.835 3.145 ;
        RECT 21.245 2.635 23.835 2.805 ;
        RECT 21.245 2.295 21.600 2.465 ;
        RECT 20.785 1.755 21.215 2.125 ;
        RECT 19.415 1.495 20.605 1.665 ;
        RECT 17.985 0.885 18.290 0.925 ;
        RECT 20.350 0.885 20.655 0.925 ;
        RECT 20.905 0.885 21.075 1.755 ;
        RECT 21.430 1.645 21.600 2.295 ;
        RECT 21.870 1.635 22.200 2.465 ;
        RECT 21.770 1.475 22.200 1.635 ;
        RECT 21.420 1.465 22.200 1.475 ;
        RECT 22.375 1.465 22.705 2.635 ;
        RECT 22.880 1.635 23.210 2.465 ;
        RECT 23.480 2.295 23.835 2.465 ;
        RECT 23.480 1.645 23.650 2.295 ;
        RECT 24.005 2.125 24.175 3.315 ;
        RECT 24.475 3.145 24.645 3.775 ;
        RECT 24.345 2.975 24.645 3.145 ;
        RECT 24.865 3.335 25.195 3.605 ;
        RECT 24.865 2.805 25.165 3.335 ;
        RECT 25.365 3.230 25.665 3.775 ;
        RECT 25.335 2.975 25.665 3.230 ;
        RECT 24.345 2.635 25.760 2.805 ;
        RECT 24.345 2.295 24.645 2.465 ;
        RECT 23.865 1.755 24.295 2.125 ;
        RECT 22.880 1.475 23.310 1.635 ;
        RECT 22.880 1.465 23.660 1.475 ;
        RECT 21.420 1.305 21.940 1.465 ;
        RECT 23.140 1.305 23.660 1.465 ;
        RECT 21.420 1.205 21.835 1.305 ;
        RECT 15.225 0.585 15.805 0.755 ;
        RECT 13.910 0.255 15.055 0.425 ;
        RECT 15.555 0.330 15.805 0.585 ;
        RECT 15.975 0.085 16.225 0.660 ;
        RECT 16.395 0.585 16.975 0.755 ;
        RECT 16.395 0.330 16.645 0.585 ;
        RECT 17.145 0.425 17.315 0.770 ;
        RECT 17.485 0.595 17.815 0.885 ;
        RECT 17.985 0.715 19.175 0.885 ;
        RECT 17.985 0.425 18.290 0.715 ;
        RECT 17.145 0.255 18.290 0.425 ;
        RECT 18.460 0.085 18.675 0.545 ;
        RECT 18.845 0.255 19.175 0.715 ;
        RECT 19.465 0.715 20.655 0.885 ;
        RECT 19.465 0.255 19.795 0.715 ;
        RECT 19.965 0.085 20.180 0.545 ;
        RECT 20.350 0.425 20.655 0.715 ;
        RECT 20.825 0.595 21.155 0.885 ;
        RECT 21.325 0.425 21.495 0.770 ;
        RECT 21.665 0.755 21.835 1.205 ;
        RECT 23.245 1.205 23.660 1.305 ;
        RECT 23.245 0.755 23.415 1.205 ;
        RECT 24.005 0.885 24.175 1.755 ;
        RECT 24.475 1.665 24.645 2.295 ;
        RECT 24.865 2.105 25.165 2.635 ;
        RECT 25.335 2.210 25.665 2.465 ;
        RECT 24.865 1.835 25.195 2.105 ;
        RECT 25.365 1.665 25.665 2.210 ;
        RECT 24.475 1.495 25.665 1.665 ;
        RECT 24.425 0.885 24.730 0.925 ;
        RECT 21.665 0.585 22.245 0.755 ;
        RECT 20.350 0.255 21.495 0.425 ;
        RECT 21.995 0.330 22.245 0.585 ;
        RECT 22.415 0.085 22.665 0.660 ;
        RECT 22.835 0.585 23.415 0.755 ;
        RECT 22.835 0.330 23.085 0.585 ;
        RECT 23.585 0.425 23.755 0.770 ;
        RECT 23.925 0.595 24.255 0.885 ;
        RECT 24.425 0.715 25.615 0.885 ;
        RECT 24.425 0.425 24.730 0.715 ;
        RECT 23.585 0.255 24.730 0.425 ;
        RECT 24.900 0.085 25.115 0.545 ;
        RECT 25.285 0.255 25.615 0.715 ;
        RECT 0.000 -0.085 25.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 5.355 0.315 5.525 ;
        RECT 0.605 5.355 0.775 5.525 ;
        RECT 1.065 5.355 1.235 5.525 ;
        RECT 1.525 5.355 1.695 5.525 ;
        RECT 1.985 5.355 2.155 5.525 ;
        RECT 2.445 5.355 2.615 5.525 ;
        RECT 2.905 5.355 3.075 5.525 ;
        RECT 3.365 5.355 3.535 5.525 ;
        RECT 3.825 5.355 3.995 5.525 ;
        RECT 4.285 5.355 4.455 5.525 ;
        RECT 4.745 5.355 4.915 5.525 ;
        RECT 5.205 5.355 5.375 5.525 ;
        RECT 5.665 5.355 5.835 5.525 ;
        RECT 6.125 5.355 6.295 5.525 ;
        RECT 6.585 5.355 6.755 5.525 ;
        RECT 7.045 5.355 7.215 5.525 ;
        RECT 7.505 5.355 7.675 5.525 ;
        RECT 7.965 5.355 8.135 5.525 ;
        RECT 8.425 5.355 8.595 5.525 ;
        RECT 8.885 5.355 9.055 5.525 ;
        RECT 9.345 5.355 9.515 5.525 ;
        RECT 9.805 5.355 9.975 5.525 ;
        RECT 10.265 5.355 10.435 5.525 ;
        RECT 10.725 5.355 10.895 5.525 ;
        RECT 11.185 5.355 11.355 5.525 ;
        RECT 11.645 5.355 11.815 5.525 ;
        RECT 12.105 5.355 12.275 5.525 ;
        RECT 12.565 5.355 12.735 5.525 ;
        RECT 13.025 5.355 13.195 5.525 ;
        RECT 13.485 5.355 13.655 5.525 ;
        RECT 13.945 5.355 14.115 5.525 ;
        RECT 14.405 5.355 14.575 5.525 ;
        RECT 14.865 5.355 15.035 5.525 ;
        RECT 15.325 5.355 15.495 5.525 ;
        RECT 15.785 5.355 15.955 5.525 ;
        RECT 16.245 5.355 16.415 5.525 ;
        RECT 16.705 5.355 16.875 5.525 ;
        RECT 17.165 5.355 17.335 5.525 ;
        RECT 17.625 5.355 17.795 5.525 ;
        RECT 18.085 5.355 18.255 5.525 ;
        RECT 18.545 5.355 18.715 5.525 ;
        RECT 19.005 5.355 19.175 5.525 ;
        RECT 19.465 5.355 19.635 5.525 ;
        RECT 19.925 5.355 20.095 5.525 ;
        RECT 20.385 5.355 20.555 5.525 ;
        RECT 20.845 5.355 21.015 5.525 ;
        RECT 21.305 5.355 21.475 5.525 ;
        RECT 21.765 5.355 21.935 5.525 ;
        RECT 22.225 5.355 22.395 5.525 ;
        RECT 22.685 5.355 22.855 5.525 ;
        RECT 23.145 5.355 23.315 5.525 ;
        RECT 23.605 5.355 23.775 5.525 ;
        RECT 24.065 5.355 24.235 5.525 ;
        RECT 24.525 5.355 24.695 5.525 ;
        RECT 24.985 5.355 25.155 5.525 ;
        RECT 25.445 5.355 25.615 5.525 ;
        RECT 0.175 3.130 0.345 3.300 ;
        RECT 1.525 3.485 1.695 3.655 ;
        RECT 1.115 3.130 1.285 3.300 ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 0.175 2.140 0.345 2.310 ;
        RECT 1.115 2.140 1.285 2.310 ;
        RECT 2.110 3.130 2.280 3.300 ;
        RECT 4.745 3.485 4.915 3.655 ;
        RECT 4.160 3.130 4.330 3.300 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 2.110 2.140 2.280 2.310 ;
        RECT 1.525 1.785 1.695 1.955 ;
        RECT 4.160 2.140 4.330 2.310 ;
        RECT 5.155 3.130 5.325 3.300 ;
        RECT 6.095 3.130 6.265 3.300 ;
        RECT 6.615 3.130 6.785 3.300 ;
        RECT 7.965 3.485 8.135 3.655 ;
        RECT 7.555 3.130 7.725 3.300 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 5.155 2.140 5.325 2.310 ;
        RECT 4.745 1.785 4.915 1.955 ;
        RECT 6.095 2.140 6.265 2.310 ;
        RECT 6.615 2.140 6.785 2.310 ;
        RECT 7.555 2.140 7.725 2.310 ;
        RECT 8.550 3.130 8.720 3.300 ;
        RECT 11.185 3.485 11.355 3.655 ;
        RECT 10.600 3.130 10.770 3.300 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 8.550 2.140 8.720 2.310 ;
        RECT 7.965 1.785 8.135 1.955 ;
        RECT 10.600 2.140 10.770 2.310 ;
        RECT 11.595 3.130 11.765 3.300 ;
        RECT 12.535 3.130 12.705 3.300 ;
        RECT 13.055 3.130 13.225 3.300 ;
        RECT 14.405 3.485 14.575 3.655 ;
        RECT 13.995 3.130 14.165 3.300 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 11.595 2.140 11.765 2.310 ;
        RECT 11.185 1.785 11.355 1.955 ;
        RECT 12.535 2.140 12.705 2.310 ;
        RECT 13.055 2.140 13.225 2.310 ;
        RECT 13.995 2.140 14.165 2.310 ;
        RECT 14.990 3.130 15.160 3.300 ;
        RECT 17.625 3.485 17.795 3.655 ;
        RECT 17.040 3.130 17.210 3.300 ;
        RECT 14.865 2.635 15.035 2.805 ;
        RECT 15.325 2.635 15.495 2.805 ;
        RECT 15.785 2.635 15.955 2.805 ;
        RECT 16.245 2.635 16.415 2.805 ;
        RECT 16.705 2.635 16.875 2.805 ;
        RECT 17.165 2.635 17.335 2.805 ;
        RECT 14.990 2.140 15.160 2.310 ;
        RECT 14.405 1.785 14.575 1.955 ;
        RECT 17.040 2.140 17.210 2.310 ;
        RECT 18.035 3.130 18.205 3.300 ;
        RECT 18.975 3.130 19.145 3.300 ;
        RECT 19.495 3.130 19.665 3.300 ;
        RECT 20.845 3.485 21.015 3.655 ;
        RECT 20.435 3.130 20.605 3.300 ;
        RECT 18.085 2.635 18.255 2.805 ;
        RECT 18.545 2.635 18.715 2.805 ;
        RECT 19.005 2.635 19.175 2.805 ;
        RECT 19.465 2.635 19.635 2.805 ;
        RECT 19.925 2.635 20.095 2.805 ;
        RECT 20.385 2.635 20.555 2.805 ;
        RECT 18.035 2.140 18.205 2.310 ;
        RECT 17.625 1.785 17.795 1.955 ;
        RECT 18.975 2.140 19.145 2.310 ;
        RECT 19.495 2.140 19.665 2.310 ;
        RECT 20.435 2.140 20.605 2.310 ;
        RECT 21.430 3.130 21.600 3.300 ;
        RECT 24.065 3.485 24.235 3.655 ;
        RECT 23.480 3.130 23.650 3.300 ;
        RECT 21.305 2.635 21.475 2.805 ;
        RECT 21.765 2.635 21.935 2.805 ;
        RECT 22.225 2.635 22.395 2.805 ;
        RECT 22.685 2.635 22.855 2.805 ;
        RECT 23.145 2.635 23.315 2.805 ;
        RECT 23.605 2.635 23.775 2.805 ;
        RECT 21.430 2.140 21.600 2.310 ;
        RECT 20.845 1.785 21.015 1.955 ;
        RECT 23.480 2.140 23.650 2.310 ;
        RECT 24.475 3.130 24.645 3.300 ;
        RECT 25.415 3.130 25.585 3.300 ;
        RECT 24.525 2.635 24.695 2.805 ;
        RECT 24.985 2.635 25.155 2.805 ;
        RECT 25.445 2.635 25.615 2.805 ;
        RECT 24.475 2.140 24.645 2.310 ;
        RECT 24.065 1.785 24.235 1.955 ;
        RECT 25.415 2.140 25.585 2.310 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
        RECT 14.405 -0.085 14.575 0.085 ;
        RECT 14.865 -0.085 15.035 0.085 ;
        RECT 15.325 -0.085 15.495 0.085 ;
        RECT 15.785 -0.085 15.955 0.085 ;
        RECT 16.245 -0.085 16.415 0.085 ;
        RECT 16.705 -0.085 16.875 0.085 ;
        RECT 17.165 -0.085 17.335 0.085 ;
        RECT 17.625 -0.085 17.795 0.085 ;
        RECT 18.085 -0.085 18.255 0.085 ;
        RECT 18.545 -0.085 18.715 0.085 ;
        RECT 19.005 -0.085 19.175 0.085 ;
        RECT 19.465 -0.085 19.635 0.085 ;
        RECT 19.925 -0.085 20.095 0.085 ;
        RECT 20.385 -0.085 20.555 0.085 ;
        RECT 20.845 -0.085 21.015 0.085 ;
        RECT 21.305 -0.085 21.475 0.085 ;
        RECT 21.765 -0.085 21.935 0.085 ;
        RECT 22.225 -0.085 22.395 0.085 ;
        RECT 22.685 -0.085 22.855 0.085 ;
        RECT 23.145 -0.085 23.315 0.085 ;
        RECT 23.605 -0.085 23.775 0.085 ;
        RECT 24.065 -0.085 24.235 0.085 ;
        RECT 24.525 -0.085 24.695 0.085 ;
        RECT 24.985 -0.085 25.155 0.085 ;
        RECT 25.445 -0.085 25.615 0.085 ;
      LAYER met1 ;
        RECT 0.115 3.285 0.405 3.330 ;
        RECT 1.055 3.285 1.345 3.330 ;
        RECT 2.050 3.285 2.340 3.330 ;
        RECT 0.115 3.145 2.340 3.285 ;
        RECT 0.115 3.100 0.405 3.145 ;
        RECT 1.055 3.100 1.345 3.145 ;
        RECT 2.050 3.100 2.340 3.145 ;
        RECT 4.100 3.285 4.390 3.330 ;
        RECT 5.095 3.285 5.385 3.330 ;
        RECT 6.035 3.285 6.325 3.330 ;
        RECT 4.100 3.145 6.325 3.285 ;
        RECT 4.100 3.100 4.390 3.145 ;
        RECT 5.095 3.100 5.385 3.145 ;
        RECT 6.035 3.100 6.325 3.145 ;
        RECT 6.555 3.285 6.845 3.330 ;
        RECT 7.495 3.285 7.785 3.330 ;
        RECT 8.490 3.285 8.780 3.330 ;
        RECT 6.555 3.145 8.780 3.285 ;
        RECT 6.555 3.100 6.845 3.145 ;
        RECT 7.495 3.100 7.785 3.145 ;
        RECT 8.490 3.100 8.780 3.145 ;
        RECT 10.540 3.285 10.830 3.330 ;
        RECT 11.535 3.285 11.825 3.330 ;
        RECT 12.475 3.285 12.765 3.330 ;
        RECT 10.540 3.145 12.765 3.285 ;
        RECT 10.540 3.100 10.830 3.145 ;
        RECT 11.535 3.100 11.825 3.145 ;
        RECT 12.475 3.100 12.765 3.145 ;
        RECT 12.995 3.285 13.285 3.330 ;
        RECT 13.935 3.285 14.225 3.330 ;
        RECT 14.930 3.285 15.220 3.330 ;
        RECT 12.995 3.145 15.220 3.285 ;
        RECT 12.995 3.100 13.285 3.145 ;
        RECT 13.935 3.100 14.225 3.145 ;
        RECT 14.930 3.100 15.220 3.145 ;
        RECT 16.980 3.285 17.270 3.330 ;
        RECT 17.975 3.285 18.265 3.330 ;
        RECT 18.915 3.285 19.205 3.330 ;
        RECT 16.980 3.145 19.205 3.285 ;
        RECT 16.980 3.100 17.270 3.145 ;
        RECT 17.975 3.100 18.265 3.145 ;
        RECT 18.915 3.100 19.205 3.145 ;
        RECT 19.435 3.285 19.725 3.330 ;
        RECT 20.375 3.285 20.665 3.330 ;
        RECT 21.370 3.285 21.660 3.330 ;
        RECT 19.435 3.145 21.660 3.285 ;
        RECT 19.435 3.100 19.725 3.145 ;
        RECT 20.375 3.100 20.665 3.145 ;
        RECT 21.370 3.100 21.660 3.145 ;
        RECT 23.420 3.285 23.710 3.330 ;
        RECT 24.415 3.285 24.705 3.330 ;
        RECT 25.355 3.285 25.645 3.330 ;
        RECT 23.420 3.145 25.645 3.285 ;
        RECT 23.420 3.100 23.710 3.145 ;
        RECT 24.415 3.100 24.705 3.145 ;
        RECT 25.355 3.100 25.645 3.145 ;
        RECT 0.115 2.295 0.405 2.340 ;
        RECT 1.055 2.295 1.345 2.340 ;
        RECT 2.050 2.295 2.340 2.340 ;
        RECT 0.115 2.155 2.340 2.295 ;
        RECT 0.115 2.110 0.405 2.155 ;
        RECT 1.055 2.110 1.345 2.155 ;
        RECT 2.050 2.110 2.340 2.155 ;
        RECT 4.100 2.295 4.390 2.340 ;
        RECT 5.095 2.295 5.385 2.340 ;
        RECT 6.035 2.295 6.325 2.340 ;
        RECT 4.100 2.155 6.325 2.295 ;
        RECT 4.100 2.110 4.390 2.155 ;
        RECT 5.095 2.110 5.385 2.155 ;
        RECT 6.035 2.110 6.325 2.155 ;
        RECT 6.555 2.295 6.845 2.340 ;
        RECT 7.495 2.295 7.785 2.340 ;
        RECT 8.490 2.295 8.780 2.340 ;
        RECT 6.555 2.155 8.780 2.295 ;
        RECT 6.555 2.110 6.845 2.155 ;
        RECT 7.495 2.110 7.785 2.155 ;
        RECT 8.490 2.110 8.780 2.155 ;
        RECT 10.540 2.295 10.830 2.340 ;
        RECT 11.535 2.295 11.825 2.340 ;
        RECT 12.475 2.295 12.765 2.340 ;
        RECT 10.540 2.155 12.765 2.295 ;
        RECT 10.540 2.110 10.830 2.155 ;
        RECT 11.535 2.110 11.825 2.155 ;
        RECT 12.475 2.110 12.765 2.155 ;
        RECT 12.995 2.295 13.285 2.340 ;
        RECT 13.935 2.295 14.225 2.340 ;
        RECT 14.930 2.295 15.220 2.340 ;
        RECT 12.995 2.155 15.220 2.295 ;
        RECT 12.995 2.110 13.285 2.155 ;
        RECT 13.935 2.110 14.225 2.155 ;
        RECT 14.930 2.110 15.220 2.155 ;
        RECT 16.980 2.295 17.270 2.340 ;
        RECT 17.975 2.295 18.265 2.340 ;
        RECT 18.915 2.295 19.205 2.340 ;
        RECT 16.980 2.155 19.205 2.295 ;
        RECT 16.980 2.110 17.270 2.155 ;
        RECT 17.975 2.110 18.265 2.155 ;
        RECT 18.915 2.110 19.205 2.155 ;
        RECT 19.435 2.295 19.725 2.340 ;
        RECT 20.375 2.295 20.665 2.340 ;
        RECT 21.370 2.295 21.660 2.340 ;
        RECT 19.435 2.155 21.660 2.295 ;
        RECT 19.435 2.110 19.725 2.155 ;
        RECT 20.375 2.110 20.665 2.155 ;
        RECT 21.370 2.110 21.660 2.155 ;
        RECT 23.420 2.295 23.710 2.340 ;
        RECT 24.415 2.295 24.705 2.340 ;
        RECT 25.355 2.295 25.645 2.340 ;
        RECT 23.420 2.155 25.645 2.295 ;
        RECT 23.420 2.110 23.710 2.155 ;
        RECT 24.415 2.110 24.705 2.155 ;
        RECT 25.355 2.110 25.645 2.155 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__muxb16to1_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__muxb16to1_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__muxb16to1_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 51.980 BY 5.440 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 50.195 4.115 51.585 4.385 ;
    END
  END D[15]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 39.495 4.115 40.885 4.385 ;
    END
  END D[14]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 37.315 4.115 38.705 4.385 ;
    END
  END D[13]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 26.615 4.115 28.005 4.385 ;
    END
  END D[12]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 23.975 4.115 25.365 4.385 ;
    END
  END D[11]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 13.275 4.115 14.665 4.385 ;
    END
  END D[10]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 11.095 4.115 12.485 4.385 ;
    END
  END D[9]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.395 4.115 1.785 4.385 ;
    END
  END D[8]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 50.195 1.055 51.585 1.325 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 39.495 1.055 40.885 1.325 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 37.315 1.055 38.705 1.325 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 26.615 1.055 28.005 1.325 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 23.975 1.055 25.365 1.325 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 13.275 1.055 14.665 1.325 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 11.095 1.055 12.485 1.325 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.395 1.055 1.785 1.325 ;
    END
  END D[0]
  PIN S[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.733200 ;
    PORT
      LAYER li1 ;
        RECT 45.625 4.115 46.220 4.445 ;
    END
  END S[15]
  PIN S[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.733200 ;
    PORT
      LAYER li1 ;
        RECT 44.860 4.115 45.455 4.445 ;
    END
  END S[14]
  PIN S[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.733200 ;
    PORT
      LAYER li1 ;
        RECT 32.745 4.115 33.340 4.445 ;
    END
  END S[13]
  PIN S[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.733200 ;
    PORT
      LAYER li1 ;
        RECT 31.980 4.115 32.575 4.445 ;
    END
  END S[12]
  PIN S[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.733200 ;
    PORT
      LAYER li1 ;
        RECT 19.405 4.115 20.000 4.445 ;
    END
  END S[11]
  PIN S[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.733200 ;
    PORT
      LAYER li1 ;
        RECT 18.640 4.115 19.235 4.445 ;
    END
  END S[10]
  PIN S[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.733200 ;
    PORT
      LAYER li1 ;
        RECT 6.525 4.115 7.120 4.445 ;
    END
  END S[9]
  PIN S[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.733200 ;
    PORT
      LAYER li1 ;
        RECT 5.760 4.115 6.355 4.445 ;
    END
  END S[8]
  PIN S[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.733200 ;
    PORT
      LAYER li1 ;
        RECT 45.625 0.995 46.220 1.325 ;
    END
  END S[7]
  PIN S[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.733200 ;
    PORT
      LAYER li1 ;
        RECT 44.860 0.995 45.455 1.325 ;
    END
  END S[6]
  PIN S[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.733200 ;
    PORT
      LAYER li1 ;
        RECT 32.745 0.995 33.340 1.325 ;
    END
  END S[5]
  PIN S[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.733200 ;
    PORT
      LAYER li1 ;
        RECT 31.980 0.995 32.575 1.325 ;
    END
  END S[4]
  PIN S[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.733200 ;
    PORT
      LAYER li1 ;
        RECT 19.405 0.995 20.000 1.325 ;
    END
  END S[3]
  PIN S[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.733200 ;
    PORT
      LAYER li1 ;
        RECT 18.640 0.995 19.235 1.325 ;
    END
  END S[2]
  PIN S[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.733200 ;
    PORT
      LAYER li1 ;
        RECT 6.525 0.995 7.120 1.325 ;
    END
  END S[1]
  PIN S[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.733200 ;
    PORT
      LAYER li1 ;
        RECT 5.760 0.995 6.355 1.325 ;
    END
  END S[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 51.980 0.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 5.200 51.980 5.680 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.980 2.345 1.015 ;
        RECT 10.535 0.980 15.225 1.015 ;
        RECT 23.415 0.980 28.565 1.015 ;
        RECT 36.755 0.980 41.445 1.015 ;
        RECT 49.635 0.980 51.975 1.015 ;
        RECT 0.005 0.785 4.545 0.980 ;
        RECT 8.335 0.785 17.425 0.980 ;
        RECT 21.215 0.785 30.765 0.980 ;
        RECT 34.555 0.785 43.645 0.980 ;
        RECT 47.435 0.785 51.975 0.980 ;
        RECT 0.005 0.200 51.975 0.785 ;
        RECT 0.005 0.105 2.345 0.200 ;
        RECT 4.910 0.105 7.970 0.200 ;
        RECT 10.535 0.105 15.225 0.200 ;
        RECT 17.790 0.105 20.850 0.200 ;
        RECT 23.415 0.105 28.565 0.200 ;
        RECT 31.130 0.105 34.190 0.200 ;
        RECT 36.755 0.105 41.445 0.200 ;
        RECT 44.010 0.105 47.070 0.200 ;
        RECT 49.635 0.105 51.975 0.200 ;
        RECT 0.145 -0.085 0.315 0.105 ;
        RECT 12.565 -0.085 13.195 0.105 ;
        RECT 25.445 -0.085 26.535 0.105 ;
        RECT 38.785 -0.085 39.415 0.105 ;
        RECT 51.665 -0.085 51.835 0.105 ;
      LAYER li1 ;
        RECT 25.845 0.265 26.135 0.810 ;
    END
    PORT
      LAYER pwell ;
        RECT 0.145 5.335 0.315 5.525 ;
        RECT 12.565 5.335 13.195 5.525 ;
        RECT 25.445 5.335 26.535 5.525 ;
        RECT 38.785 5.335 39.415 5.525 ;
        RECT 51.665 5.335 51.835 5.525 ;
        RECT 0.005 5.240 2.345 5.335 ;
        RECT 4.910 5.240 7.970 5.335 ;
        RECT 10.535 5.240 15.225 5.335 ;
        RECT 17.790 5.240 20.850 5.335 ;
        RECT 23.415 5.240 28.565 5.335 ;
        RECT 31.130 5.240 34.190 5.335 ;
        RECT 36.755 5.240 41.445 5.335 ;
        RECT 44.010 5.240 47.070 5.335 ;
        RECT 49.635 5.240 51.975 5.335 ;
        RECT 0.005 4.655 51.975 5.240 ;
        RECT 0.005 4.460 4.545 4.655 ;
        RECT 8.335 4.460 17.425 4.655 ;
        RECT 21.215 4.460 30.765 4.655 ;
        RECT 34.555 4.460 43.645 4.655 ;
        RECT 47.435 4.460 51.975 4.655 ;
        RECT 0.005 4.425 2.345 4.460 ;
        RECT 10.535 4.425 15.225 4.460 ;
        RECT 23.415 4.425 28.565 4.460 ;
        RECT 36.755 4.425 41.445 4.460 ;
        RECT 49.635 4.425 51.975 4.460 ;
      LAYER li1 ;
        RECT 25.845 4.630 26.135 5.175 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 52.170 4.135 ;
      LAYER li1 ;
        RECT 25.845 2.985 26.135 3.970 ;
        RECT 25.845 1.470 26.135 2.455 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 51.980 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.102400 ;
    PORT
      LAYER met1 ;
        RECT 2.985 3.640 3.275 3.685 ;
        RECT 3.925 3.640 4.215 3.685 ;
        RECT 8.665 3.640 8.955 3.685 ;
        RECT 9.605 3.640 9.895 3.685 ;
        RECT 15.865 3.640 16.155 3.685 ;
        RECT 16.805 3.640 17.095 3.685 ;
        RECT 21.545 3.640 21.835 3.685 ;
        RECT 22.485 3.640 22.775 3.685 ;
        RECT 29.205 3.640 29.495 3.685 ;
        RECT 30.145 3.640 30.435 3.685 ;
        RECT 34.885 3.640 35.175 3.685 ;
        RECT 35.825 3.640 36.115 3.685 ;
        RECT 42.085 3.640 42.375 3.685 ;
        RECT 43.025 3.640 43.315 3.685 ;
        RECT 47.765 3.640 48.055 3.685 ;
        RECT 48.705 3.640 48.995 3.685 ;
        RECT 2.985 3.500 48.995 3.640 ;
        RECT 2.985 3.455 3.275 3.500 ;
        RECT 3.925 3.455 4.215 3.500 ;
        RECT 8.665 3.455 8.955 3.500 ;
        RECT 9.605 3.455 9.895 3.500 ;
        RECT 15.865 3.455 16.155 3.500 ;
        RECT 16.805 3.455 17.095 3.500 ;
        RECT 21.545 3.455 21.835 3.500 ;
        RECT 22.485 3.455 22.775 3.500 ;
        RECT 29.205 3.455 29.495 3.500 ;
        RECT 30.145 3.455 30.435 3.500 ;
        RECT 34.885 3.455 35.175 3.500 ;
        RECT 35.825 3.455 36.115 3.500 ;
        RECT 42.085 3.455 42.375 3.500 ;
        RECT 43.025 3.455 43.315 3.500 ;
        RECT 47.765 3.455 48.055 3.500 ;
        RECT 48.705 3.455 48.995 3.500 ;
        RECT 2.985 1.940 3.275 1.985 ;
        RECT 3.925 1.940 4.215 1.985 ;
        RECT 8.665 1.940 8.955 1.985 ;
        RECT 9.605 1.940 9.895 1.985 ;
        RECT 15.865 1.940 16.155 1.985 ;
        RECT 16.805 1.940 17.095 1.985 ;
        RECT 21.545 1.940 21.835 1.985 ;
        RECT 22.485 1.940 22.775 1.985 ;
        RECT 29.205 1.940 29.495 1.985 ;
        RECT 30.145 1.940 30.435 1.985 ;
        RECT 34.885 1.940 35.175 1.985 ;
        RECT 35.825 1.940 36.115 1.985 ;
        RECT 42.085 1.940 42.375 1.985 ;
        RECT 43.025 1.940 43.315 1.985 ;
        RECT 47.765 1.940 48.055 1.985 ;
        RECT 48.705 1.940 48.995 1.985 ;
        RECT 2.985 1.800 48.995 1.940 ;
        RECT 2.985 1.755 3.275 1.800 ;
        RECT 3.925 1.755 4.215 1.800 ;
        RECT 8.665 1.755 8.955 1.800 ;
        RECT 9.605 1.755 9.895 1.800 ;
        RECT 15.865 1.755 16.155 1.800 ;
        RECT 16.805 1.755 17.095 1.800 ;
        RECT 21.545 1.755 21.835 1.800 ;
        RECT 22.485 1.755 22.775 1.800 ;
        RECT 29.205 1.755 29.495 1.800 ;
        RECT 30.145 1.755 30.435 1.800 ;
        RECT 34.885 1.755 35.175 1.800 ;
        RECT 35.825 1.755 36.115 1.800 ;
        RECT 42.085 1.755 42.375 1.800 ;
        RECT 43.025 1.755 43.315 1.800 ;
        RECT 47.765 1.755 48.055 1.800 ;
        RECT 48.705 1.755 48.995 1.800 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 5.355 51.980 5.525 ;
        RECT 0.145 4.555 0.395 5.355 ;
        RECT 0.565 4.725 0.895 5.185 ;
        RECT 1.065 4.895 1.335 5.355 ;
        RECT 1.505 4.725 1.835 5.185 ;
        RECT 2.005 4.895 2.255 5.355 ;
        RECT 2.425 5.015 4.455 5.185 ;
        RECT 2.425 4.725 2.695 5.015 ;
        RECT 0.565 4.555 2.695 4.725 ;
        RECT 2.865 4.555 3.195 4.845 ;
        RECT 3.365 4.670 3.535 5.015 ;
        RECT 2.965 4.375 3.195 4.555 ;
        RECT 3.705 4.375 4.035 4.845 ;
        RECT 4.205 4.670 4.455 5.015 ;
        RECT 4.960 4.830 5.250 5.355 ;
        RECT 5.420 4.615 5.670 5.160 ;
        RECT 5.880 4.830 6.170 5.355 ;
        RECT 6.710 4.830 7.000 5.355 ;
        RECT 7.210 4.615 7.460 5.160 ;
        RECT 7.630 4.830 7.920 5.355 ;
        RECT 8.425 5.015 10.455 5.185 ;
        RECT 8.425 4.670 8.675 5.015 ;
        RECT 5.420 4.375 5.590 4.615 ;
        RECT 2.965 4.075 4.235 4.375 ;
        RECT 0.125 2.805 0.395 3.945 ;
        RECT 0.565 3.775 2.795 3.945 ;
        RECT 0.565 2.975 0.895 3.775 ;
        RECT 1.065 2.805 1.335 3.605 ;
        RECT 1.505 2.975 1.835 3.775 ;
        RECT 2.005 2.805 2.275 3.605 ;
        RECT 2.495 2.975 2.795 3.775 ;
        RECT 0.000 2.635 2.795 2.805 ;
        RECT 0.125 1.495 0.395 2.635 ;
        RECT 0.565 1.665 0.895 2.465 ;
        RECT 1.065 1.835 1.335 2.635 ;
        RECT 1.505 1.665 1.835 2.465 ;
        RECT 2.005 1.835 2.275 2.635 ;
        RECT 2.495 1.665 2.795 2.465 ;
        RECT 0.565 1.495 2.795 1.665 ;
        RECT 2.965 1.365 3.295 4.075 ;
        RECT 3.465 2.975 3.735 3.905 ;
        RECT 3.465 1.535 3.735 2.465 ;
        RECT 3.905 1.365 4.235 4.075 ;
        RECT 4.405 4.045 5.590 4.375 ;
        RECT 4.405 2.975 4.705 3.875 ;
        RECT 5.420 3.835 5.590 4.045 ;
        RECT 7.290 4.375 7.460 4.615 ;
        RECT 8.845 4.375 9.175 4.845 ;
        RECT 9.345 4.670 9.515 5.015 ;
        RECT 9.685 4.555 10.015 4.845 ;
        RECT 10.185 4.725 10.455 5.015 ;
        RECT 10.625 4.895 10.875 5.355 ;
        RECT 11.045 4.725 11.375 5.185 ;
        RECT 11.545 4.895 11.815 5.355 ;
        RECT 11.985 4.725 12.315 5.185 ;
        RECT 10.185 4.555 12.315 4.725 ;
        RECT 12.485 4.555 12.735 5.355 ;
        RECT 13.025 4.555 13.275 5.355 ;
        RECT 13.445 4.725 13.775 5.185 ;
        RECT 13.945 4.895 14.215 5.355 ;
        RECT 14.385 4.725 14.715 5.185 ;
        RECT 14.885 4.895 15.135 5.355 ;
        RECT 15.305 5.015 17.335 5.185 ;
        RECT 15.305 4.725 15.575 5.015 ;
        RECT 13.445 4.555 15.575 4.725 ;
        RECT 15.745 4.555 16.075 4.845 ;
        RECT 16.245 4.670 16.415 5.015 ;
        RECT 9.685 4.375 9.915 4.555 ;
        RECT 7.290 4.045 8.475 4.375 ;
        RECT 8.645 4.075 9.915 4.375 ;
        RECT 7.290 3.835 7.460 4.045 ;
        RECT 4.950 2.805 5.225 3.835 ;
        RECT 5.420 2.975 5.750 3.835 ;
        RECT 5.920 2.805 6.220 3.835 ;
        RECT 6.660 2.805 6.960 3.835 ;
        RECT 7.130 2.975 7.460 3.835 ;
        RECT 7.655 2.805 7.930 3.835 ;
        RECT 8.175 2.975 8.475 3.875 ;
        RECT 4.405 2.635 8.475 2.805 ;
        RECT 4.405 1.565 4.705 2.465 ;
        RECT 4.950 1.605 5.225 2.635 ;
        RECT 5.420 1.605 5.750 2.465 ;
        RECT 5.920 1.605 6.220 2.635 ;
        RECT 6.660 1.605 6.960 2.635 ;
        RECT 7.130 1.605 7.460 2.465 ;
        RECT 7.655 1.605 7.930 2.635 ;
        RECT 5.420 1.395 5.590 1.605 ;
        RECT 2.965 1.065 4.235 1.365 ;
        RECT 4.405 1.065 5.590 1.395 ;
        RECT 2.965 0.885 3.195 1.065 ;
        RECT 0.145 0.085 0.395 0.885 ;
        RECT 0.565 0.715 2.695 0.885 ;
        RECT 0.565 0.255 0.895 0.715 ;
        RECT 1.065 0.085 1.335 0.545 ;
        RECT 1.505 0.255 1.835 0.715 ;
        RECT 2.005 0.085 2.255 0.545 ;
        RECT 2.425 0.425 2.695 0.715 ;
        RECT 2.865 0.595 3.195 0.885 ;
        RECT 3.365 0.425 3.535 0.770 ;
        RECT 3.705 0.595 4.035 1.065 ;
        RECT 5.420 0.825 5.590 1.065 ;
        RECT 7.290 1.395 7.460 1.605 ;
        RECT 8.175 1.565 8.475 2.465 ;
        RECT 7.290 1.065 8.475 1.395 ;
        RECT 8.645 1.365 8.975 4.075 ;
        RECT 9.145 2.975 9.415 3.905 ;
        RECT 9.145 1.535 9.415 2.465 ;
        RECT 9.585 1.365 9.915 4.075 ;
        RECT 15.845 4.375 16.075 4.555 ;
        RECT 16.585 4.375 16.915 4.845 ;
        RECT 17.085 4.670 17.335 5.015 ;
        RECT 17.840 4.830 18.130 5.355 ;
        RECT 18.300 4.615 18.550 5.160 ;
        RECT 18.760 4.830 19.050 5.355 ;
        RECT 19.590 4.830 19.880 5.355 ;
        RECT 20.090 4.615 20.340 5.160 ;
        RECT 20.510 4.830 20.800 5.355 ;
        RECT 21.305 5.015 23.335 5.185 ;
        RECT 21.305 4.670 21.555 5.015 ;
        RECT 18.300 4.375 18.470 4.615 ;
        RECT 15.845 4.075 17.115 4.375 ;
        RECT 10.085 3.775 12.315 3.945 ;
        RECT 10.085 2.975 10.385 3.775 ;
        RECT 10.605 2.805 10.875 3.605 ;
        RECT 11.045 2.975 11.375 3.775 ;
        RECT 11.545 2.805 11.815 3.605 ;
        RECT 11.985 2.975 12.315 3.775 ;
        RECT 12.485 2.805 12.755 3.945 ;
        RECT 13.005 2.805 13.275 3.945 ;
        RECT 13.445 3.775 15.675 3.945 ;
        RECT 13.445 2.975 13.775 3.775 ;
        RECT 13.945 2.805 14.215 3.605 ;
        RECT 14.385 2.975 14.715 3.775 ;
        RECT 14.885 2.805 15.155 3.605 ;
        RECT 15.375 2.975 15.675 3.775 ;
        RECT 10.085 2.635 15.675 2.805 ;
        RECT 10.085 1.665 10.385 2.465 ;
        RECT 10.605 1.835 10.875 2.635 ;
        RECT 11.045 1.665 11.375 2.465 ;
        RECT 11.545 1.835 11.815 2.635 ;
        RECT 11.985 1.665 12.315 2.465 ;
        RECT 10.085 1.495 12.315 1.665 ;
        RECT 12.485 1.495 12.755 2.635 ;
        RECT 13.005 1.495 13.275 2.635 ;
        RECT 13.445 1.665 13.775 2.465 ;
        RECT 13.945 1.835 14.215 2.635 ;
        RECT 14.385 1.665 14.715 2.465 ;
        RECT 14.885 1.835 15.155 2.635 ;
        RECT 15.375 1.665 15.675 2.465 ;
        RECT 13.445 1.495 15.675 1.665 ;
        RECT 8.645 1.065 9.915 1.365 ;
        RECT 7.290 0.825 7.460 1.065 ;
        RECT 4.205 0.425 4.455 0.770 ;
        RECT 2.425 0.255 4.455 0.425 ;
        RECT 4.960 0.085 5.250 0.610 ;
        RECT 5.420 0.280 5.670 0.825 ;
        RECT 5.880 0.085 6.170 0.610 ;
        RECT 6.710 0.085 7.000 0.610 ;
        RECT 7.210 0.280 7.460 0.825 ;
        RECT 7.630 0.085 7.920 0.610 ;
        RECT 8.425 0.425 8.675 0.770 ;
        RECT 8.845 0.595 9.175 1.065 ;
        RECT 9.685 0.885 9.915 1.065 ;
        RECT 15.845 1.365 16.175 4.075 ;
        RECT 16.345 2.975 16.615 3.905 ;
        RECT 16.345 1.535 16.615 2.465 ;
        RECT 16.785 1.365 17.115 4.075 ;
        RECT 17.285 4.045 18.470 4.375 ;
        RECT 17.285 2.975 17.585 3.875 ;
        RECT 18.300 3.835 18.470 4.045 ;
        RECT 20.170 4.375 20.340 4.615 ;
        RECT 21.725 4.375 22.055 4.845 ;
        RECT 22.225 4.670 22.395 5.015 ;
        RECT 22.565 4.555 22.895 4.845 ;
        RECT 23.065 4.725 23.335 5.015 ;
        RECT 23.505 4.895 23.755 5.355 ;
        RECT 23.925 4.725 24.255 5.185 ;
        RECT 24.425 4.895 24.695 5.355 ;
        RECT 24.865 4.725 25.195 5.185 ;
        RECT 23.065 4.555 25.195 4.725 ;
        RECT 25.365 4.555 25.615 5.355 ;
        RECT 26.365 4.555 26.615 5.355 ;
        RECT 26.785 4.725 27.115 5.185 ;
        RECT 27.285 4.895 27.555 5.355 ;
        RECT 27.725 4.725 28.055 5.185 ;
        RECT 28.225 4.895 28.475 5.355 ;
        RECT 28.645 5.015 30.675 5.185 ;
        RECT 28.645 4.725 28.915 5.015 ;
        RECT 26.785 4.555 28.915 4.725 ;
        RECT 29.085 4.555 29.415 4.845 ;
        RECT 29.585 4.670 29.755 5.015 ;
        RECT 22.565 4.375 22.795 4.555 ;
        RECT 20.170 4.045 21.355 4.375 ;
        RECT 21.525 4.075 22.795 4.375 ;
        RECT 20.170 3.835 20.340 4.045 ;
        RECT 17.830 2.805 18.105 3.835 ;
        RECT 18.300 2.975 18.630 3.835 ;
        RECT 18.800 2.805 19.100 3.835 ;
        RECT 19.540 2.805 19.840 3.835 ;
        RECT 20.010 2.975 20.340 3.835 ;
        RECT 20.535 2.805 20.810 3.835 ;
        RECT 21.055 2.975 21.355 3.875 ;
        RECT 17.285 2.635 21.355 2.805 ;
        RECT 17.285 1.565 17.585 2.465 ;
        RECT 17.830 1.605 18.105 2.635 ;
        RECT 18.300 1.605 18.630 2.465 ;
        RECT 18.800 1.605 19.100 2.635 ;
        RECT 19.540 1.605 19.840 2.635 ;
        RECT 20.010 1.605 20.340 2.465 ;
        RECT 20.535 1.605 20.810 2.635 ;
        RECT 18.300 1.395 18.470 1.605 ;
        RECT 15.845 1.065 17.115 1.365 ;
        RECT 17.285 1.065 18.470 1.395 ;
        RECT 15.845 0.885 16.075 1.065 ;
        RECT 9.345 0.425 9.515 0.770 ;
        RECT 9.685 0.595 10.015 0.885 ;
        RECT 10.185 0.715 12.315 0.885 ;
        RECT 10.185 0.425 10.455 0.715 ;
        RECT 8.425 0.255 10.455 0.425 ;
        RECT 10.625 0.085 10.875 0.545 ;
        RECT 11.045 0.255 11.375 0.715 ;
        RECT 11.545 0.085 11.815 0.545 ;
        RECT 11.985 0.255 12.315 0.715 ;
        RECT 12.485 0.085 12.735 0.885 ;
        RECT 13.025 0.085 13.275 0.885 ;
        RECT 13.445 0.715 15.575 0.885 ;
        RECT 13.445 0.255 13.775 0.715 ;
        RECT 13.945 0.085 14.215 0.545 ;
        RECT 14.385 0.255 14.715 0.715 ;
        RECT 14.885 0.085 15.135 0.545 ;
        RECT 15.305 0.425 15.575 0.715 ;
        RECT 15.745 0.595 16.075 0.885 ;
        RECT 16.245 0.425 16.415 0.770 ;
        RECT 16.585 0.595 16.915 1.065 ;
        RECT 18.300 0.825 18.470 1.065 ;
        RECT 20.170 1.395 20.340 1.605 ;
        RECT 21.055 1.565 21.355 2.465 ;
        RECT 20.170 1.065 21.355 1.395 ;
        RECT 21.525 1.365 21.855 4.075 ;
        RECT 22.025 2.975 22.295 3.905 ;
        RECT 22.025 1.535 22.295 2.465 ;
        RECT 22.465 1.365 22.795 4.075 ;
        RECT 29.185 4.375 29.415 4.555 ;
        RECT 29.925 4.375 30.255 4.845 ;
        RECT 30.425 4.670 30.675 5.015 ;
        RECT 31.180 4.830 31.470 5.355 ;
        RECT 31.640 4.615 31.890 5.160 ;
        RECT 32.100 4.830 32.390 5.355 ;
        RECT 32.930 4.830 33.220 5.355 ;
        RECT 33.430 4.615 33.680 5.160 ;
        RECT 33.850 4.830 34.140 5.355 ;
        RECT 34.645 5.015 36.675 5.185 ;
        RECT 34.645 4.670 34.895 5.015 ;
        RECT 31.640 4.375 31.810 4.615 ;
        RECT 29.185 4.075 30.455 4.375 ;
        RECT 22.965 3.775 25.195 3.945 ;
        RECT 22.965 2.975 23.265 3.775 ;
        RECT 23.485 2.805 23.755 3.605 ;
        RECT 23.925 2.975 24.255 3.775 ;
        RECT 24.425 2.805 24.695 3.605 ;
        RECT 24.865 2.975 25.195 3.775 ;
        RECT 25.365 2.805 25.635 3.945 ;
        RECT 26.345 2.805 26.615 3.945 ;
        RECT 26.785 3.775 29.015 3.945 ;
        RECT 26.785 2.975 27.115 3.775 ;
        RECT 27.285 2.805 27.555 3.605 ;
        RECT 27.725 2.975 28.055 3.775 ;
        RECT 28.225 2.805 28.495 3.605 ;
        RECT 28.715 2.975 29.015 3.775 ;
        RECT 22.965 2.635 29.015 2.805 ;
        RECT 22.965 1.665 23.265 2.465 ;
        RECT 23.485 1.835 23.755 2.635 ;
        RECT 23.925 1.665 24.255 2.465 ;
        RECT 24.425 1.835 24.695 2.635 ;
        RECT 24.865 1.665 25.195 2.465 ;
        RECT 22.965 1.495 25.195 1.665 ;
        RECT 25.365 1.495 25.635 2.635 ;
        RECT 26.345 1.495 26.615 2.635 ;
        RECT 26.785 1.665 27.115 2.465 ;
        RECT 27.285 1.835 27.555 2.635 ;
        RECT 27.725 1.665 28.055 2.465 ;
        RECT 28.225 1.835 28.495 2.635 ;
        RECT 28.715 1.665 29.015 2.465 ;
        RECT 26.785 1.495 29.015 1.665 ;
        RECT 21.525 1.065 22.795 1.365 ;
        RECT 20.170 0.825 20.340 1.065 ;
        RECT 17.085 0.425 17.335 0.770 ;
        RECT 15.305 0.255 17.335 0.425 ;
        RECT 17.840 0.085 18.130 0.610 ;
        RECT 18.300 0.280 18.550 0.825 ;
        RECT 18.760 0.085 19.050 0.610 ;
        RECT 19.590 0.085 19.880 0.610 ;
        RECT 20.090 0.280 20.340 0.825 ;
        RECT 20.510 0.085 20.800 0.610 ;
        RECT 21.305 0.425 21.555 0.770 ;
        RECT 21.725 0.595 22.055 1.065 ;
        RECT 22.565 0.885 22.795 1.065 ;
        RECT 29.185 1.365 29.515 4.075 ;
        RECT 29.685 2.975 29.955 3.905 ;
        RECT 29.685 1.535 29.955 2.465 ;
        RECT 30.125 1.365 30.455 4.075 ;
        RECT 30.625 4.045 31.810 4.375 ;
        RECT 30.625 2.975 30.925 3.875 ;
        RECT 31.640 3.835 31.810 4.045 ;
        RECT 33.510 4.375 33.680 4.615 ;
        RECT 35.065 4.375 35.395 4.845 ;
        RECT 35.565 4.670 35.735 5.015 ;
        RECT 35.905 4.555 36.235 4.845 ;
        RECT 36.405 4.725 36.675 5.015 ;
        RECT 36.845 4.895 37.095 5.355 ;
        RECT 37.265 4.725 37.595 5.185 ;
        RECT 37.765 4.895 38.035 5.355 ;
        RECT 38.205 4.725 38.535 5.185 ;
        RECT 36.405 4.555 38.535 4.725 ;
        RECT 38.705 4.555 38.955 5.355 ;
        RECT 39.245 4.555 39.495 5.355 ;
        RECT 39.665 4.725 39.995 5.185 ;
        RECT 40.165 4.895 40.435 5.355 ;
        RECT 40.605 4.725 40.935 5.185 ;
        RECT 41.105 4.895 41.355 5.355 ;
        RECT 41.525 5.015 43.555 5.185 ;
        RECT 41.525 4.725 41.795 5.015 ;
        RECT 39.665 4.555 41.795 4.725 ;
        RECT 41.965 4.555 42.295 4.845 ;
        RECT 42.465 4.670 42.635 5.015 ;
        RECT 35.905 4.375 36.135 4.555 ;
        RECT 33.510 4.045 34.695 4.375 ;
        RECT 34.865 4.075 36.135 4.375 ;
        RECT 33.510 3.835 33.680 4.045 ;
        RECT 31.170 2.805 31.445 3.835 ;
        RECT 31.640 2.975 31.970 3.835 ;
        RECT 32.140 2.805 32.440 3.835 ;
        RECT 32.880 2.805 33.180 3.835 ;
        RECT 33.350 2.975 33.680 3.835 ;
        RECT 33.875 2.805 34.150 3.835 ;
        RECT 34.395 2.975 34.695 3.875 ;
        RECT 30.625 2.635 34.695 2.805 ;
        RECT 30.625 1.565 30.925 2.465 ;
        RECT 31.170 1.605 31.445 2.635 ;
        RECT 31.640 1.605 31.970 2.465 ;
        RECT 32.140 1.605 32.440 2.635 ;
        RECT 32.880 1.605 33.180 2.635 ;
        RECT 33.350 1.605 33.680 2.465 ;
        RECT 33.875 1.605 34.150 2.635 ;
        RECT 31.640 1.395 31.810 1.605 ;
        RECT 29.185 1.065 30.455 1.365 ;
        RECT 30.625 1.065 31.810 1.395 ;
        RECT 29.185 0.885 29.415 1.065 ;
        RECT 22.225 0.425 22.395 0.770 ;
        RECT 22.565 0.595 22.895 0.885 ;
        RECT 23.065 0.715 25.195 0.885 ;
        RECT 23.065 0.425 23.335 0.715 ;
        RECT 21.305 0.255 23.335 0.425 ;
        RECT 23.505 0.085 23.755 0.545 ;
        RECT 23.925 0.255 24.255 0.715 ;
        RECT 24.425 0.085 24.695 0.545 ;
        RECT 24.865 0.255 25.195 0.715 ;
        RECT 25.365 0.085 25.615 0.885 ;
        RECT 26.365 0.085 26.615 0.885 ;
        RECT 26.785 0.715 28.915 0.885 ;
        RECT 26.785 0.255 27.115 0.715 ;
        RECT 27.285 0.085 27.555 0.545 ;
        RECT 27.725 0.255 28.055 0.715 ;
        RECT 28.225 0.085 28.475 0.545 ;
        RECT 28.645 0.425 28.915 0.715 ;
        RECT 29.085 0.595 29.415 0.885 ;
        RECT 29.585 0.425 29.755 0.770 ;
        RECT 29.925 0.595 30.255 1.065 ;
        RECT 31.640 0.825 31.810 1.065 ;
        RECT 33.510 1.395 33.680 1.605 ;
        RECT 34.395 1.565 34.695 2.465 ;
        RECT 33.510 1.065 34.695 1.395 ;
        RECT 34.865 1.365 35.195 4.075 ;
        RECT 35.365 2.975 35.635 3.905 ;
        RECT 35.365 1.535 35.635 2.465 ;
        RECT 35.805 1.365 36.135 4.075 ;
        RECT 42.065 4.375 42.295 4.555 ;
        RECT 42.805 4.375 43.135 4.845 ;
        RECT 43.305 4.670 43.555 5.015 ;
        RECT 44.060 4.830 44.350 5.355 ;
        RECT 44.520 4.615 44.770 5.160 ;
        RECT 44.980 4.830 45.270 5.355 ;
        RECT 45.810 4.830 46.100 5.355 ;
        RECT 46.310 4.615 46.560 5.160 ;
        RECT 46.730 4.830 47.020 5.355 ;
        RECT 47.525 5.015 49.555 5.185 ;
        RECT 47.525 4.670 47.775 5.015 ;
        RECT 44.520 4.375 44.690 4.615 ;
        RECT 42.065 4.075 43.335 4.375 ;
        RECT 36.305 3.775 38.535 3.945 ;
        RECT 36.305 2.975 36.605 3.775 ;
        RECT 36.825 2.805 37.095 3.605 ;
        RECT 37.265 2.975 37.595 3.775 ;
        RECT 37.765 2.805 38.035 3.605 ;
        RECT 38.205 2.975 38.535 3.775 ;
        RECT 38.705 2.805 38.975 3.945 ;
        RECT 39.225 2.805 39.495 3.945 ;
        RECT 39.665 3.775 41.895 3.945 ;
        RECT 39.665 2.975 39.995 3.775 ;
        RECT 40.165 2.805 40.435 3.605 ;
        RECT 40.605 2.975 40.935 3.775 ;
        RECT 41.105 2.805 41.375 3.605 ;
        RECT 41.595 2.975 41.895 3.775 ;
        RECT 36.305 2.635 41.895 2.805 ;
        RECT 36.305 1.665 36.605 2.465 ;
        RECT 36.825 1.835 37.095 2.635 ;
        RECT 37.265 1.665 37.595 2.465 ;
        RECT 37.765 1.835 38.035 2.635 ;
        RECT 38.205 1.665 38.535 2.465 ;
        RECT 36.305 1.495 38.535 1.665 ;
        RECT 38.705 1.495 38.975 2.635 ;
        RECT 39.225 1.495 39.495 2.635 ;
        RECT 39.665 1.665 39.995 2.465 ;
        RECT 40.165 1.835 40.435 2.635 ;
        RECT 40.605 1.665 40.935 2.465 ;
        RECT 41.105 1.835 41.375 2.635 ;
        RECT 41.595 1.665 41.895 2.465 ;
        RECT 39.665 1.495 41.895 1.665 ;
        RECT 34.865 1.065 36.135 1.365 ;
        RECT 33.510 0.825 33.680 1.065 ;
        RECT 30.425 0.425 30.675 0.770 ;
        RECT 28.645 0.255 30.675 0.425 ;
        RECT 31.180 0.085 31.470 0.610 ;
        RECT 31.640 0.280 31.890 0.825 ;
        RECT 32.100 0.085 32.390 0.610 ;
        RECT 32.930 0.085 33.220 0.610 ;
        RECT 33.430 0.280 33.680 0.825 ;
        RECT 33.850 0.085 34.140 0.610 ;
        RECT 34.645 0.425 34.895 0.770 ;
        RECT 35.065 0.595 35.395 1.065 ;
        RECT 35.905 0.885 36.135 1.065 ;
        RECT 42.065 1.365 42.395 4.075 ;
        RECT 42.565 2.975 42.835 3.905 ;
        RECT 42.565 1.535 42.835 2.465 ;
        RECT 43.005 1.365 43.335 4.075 ;
        RECT 43.505 4.045 44.690 4.375 ;
        RECT 43.505 2.975 43.805 3.875 ;
        RECT 44.520 3.835 44.690 4.045 ;
        RECT 46.390 4.375 46.560 4.615 ;
        RECT 47.945 4.375 48.275 4.845 ;
        RECT 48.445 4.670 48.615 5.015 ;
        RECT 48.785 4.555 49.115 4.845 ;
        RECT 49.285 4.725 49.555 5.015 ;
        RECT 49.725 4.895 49.975 5.355 ;
        RECT 50.145 4.725 50.475 5.185 ;
        RECT 50.645 4.895 50.915 5.355 ;
        RECT 51.085 4.725 51.415 5.185 ;
        RECT 49.285 4.555 51.415 4.725 ;
        RECT 51.585 4.555 51.835 5.355 ;
        RECT 48.785 4.375 49.015 4.555 ;
        RECT 46.390 4.045 47.575 4.375 ;
        RECT 47.745 4.075 49.015 4.375 ;
        RECT 46.390 3.835 46.560 4.045 ;
        RECT 44.050 2.805 44.325 3.835 ;
        RECT 44.520 2.975 44.850 3.835 ;
        RECT 45.020 2.805 45.320 3.835 ;
        RECT 45.760 2.805 46.060 3.835 ;
        RECT 46.230 2.975 46.560 3.835 ;
        RECT 46.755 2.805 47.030 3.835 ;
        RECT 47.275 2.975 47.575 3.875 ;
        RECT 43.505 2.635 47.575 2.805 ;
        RECT 43.505 1.565 43.805 2.465 ;
        RECT 44.050 1.605 44.325 2.635 ;
        RECT 44.520 1.605 44.850 2.465 ;
        RECT 45.020 1.605 45.320 2.635 ;
        RECT 45.760 1.605 46.060 2.635 ;
        RECT 46.230 1.605 46.560 2.465 ;
        RECT 46.755 1.605 47.030 2.635 ;
        RECT 44.520 1.395 44.690 1.605 ;
        RECT 42.065 1.065 43.335 1.365 ;
        RECT 43.505 1.065 44.690 1.395 ;
        RECT 42.065 0.885 42.295 1.065 ;
        RECT 35.565 0.425 35.735 0.770 ;
        RECT 35.905 0.595 36.235 0.885 ;
        RECT 36.405 0.715 38.535 0.885 ;
        RECT 36.405 0.425 36.675 0.715 ;
        RECT 34.645 0.255 36.675 0.425 ;
        RECT 36.845 0.085 37.095 0.545 ;
        RECT 37.265 0.255 37.595 0.715 ;
        RECT 37.765 0.085 38.035 0.545 ;
        RECT 38.205 0.255 38.535 0.715 ;
        RECT 38.705 0.085 38.955 0.885 ;
        RECT 39.245 0.085 39.495 0.885 ;
        RECT 39.665 0.715 41.795 0.885 ;
        RECT 39.665 0.255 39.995 0.715 ;
        RECT 40.165 0.085 40.435 0.545 ;
        RECT 40.605 0.255 40.935 0.715 ;
        RECT 41.105 0.085 41.355 0.545 ;
        RECT 41.525 0.425 41.795 0.715 ;
        RECT 41.965 0.595 42.295 0.885 ;
        RECT 42.465 0.425 42.635 0.770 ;
        RECT 42.805 0.595 43.135 1.065 ;
        RECT 44.520 0.825 44.690 1.065 ;
        RECT 46.390 1.395 46.560 1.605 ;
        RECT 47.275 1.565 47.575 2.465 ;
        RECT 46.390 1.065 47.575 1.395 ;
        RECT 47.745 1.365 48.075 4.075 ;
        RECT 48.245 2.975 48.515 3.905 ;
        RECT 48.245 1.535 48.515 2.465 ;
        RECT 48.685 1.365 49.015 4.075 ;
        RECT 49.185 3.775 51.415 3.945 ;
        RECT 49.185 2.975 49.485 3.775 ;
        RECT 49.705 2.805 49.975 3.605 ;
        RECT 50.145 2.975 50.475 3.775 ;
        RECT 50.645 2.805 50.915 3.605 ;
        RECT 51.085 2.975 51.415 3.775 ;
        RECT 51.585 2.805 51.855 3.945 ;
        RECT 49.185 2.635 51.980 2.805 ;
        RECT 49.185 1.665 49.485 2.465 ;
        RECT 49.705 1.835 49.975 2.635 ;
        RECT 50.145 1.665 50.475 2.465 ;
        RECT 50.645 1.835 50.915 2.635 ;
        RECT 51.085 1.665 51.415 2.465 ;
        RECT 49.185 1.495 51.415 1.665 ;
        RECT 51.585 1.495 51.855 2.635 ;
        RECT 47.745 1.065 49.015 1.365 ;
        RECT 46.390 0.825 46.560 1.065 ;
        RECT 43.305 0.425 43.555 0.770 ;
        RECT 41.525 0.255 43.555 0.425 ;
        RECT 44.060 0.085 44.350 0.610 ;
        RECT 44.520 0.280 44.770 0.825 ;
        RECT 44.980 0.085 45.270 0.610 ;
        RECT 45.810 0.085 46.100 0.610 ;
        RECT 46.310 0.280 46.560 0.825 ;
        RECT 46.730 0.085 47.020 0.610 ;
        RECT 47.525 0.425 47.775 0.770 ;
        RECT 47.945 0.595 48.275 1.065 ;
        RECT 48.785 0.885 49.015 1.065 ;
        RECT 48.445 0.425 48.615 0.770 ;
        RECT 48.785 0.595 49.115 0.885 ;
        RECT 49.285 0.715 51.415 0.885 ;
        RECT 49.285 0.425 49.555 0.715 ;
        RECT 47.525 0.255 49.555 0.425 ;
        RECT 49.725 0.085 49.975 0.545 ;
        RECT 50.145 0.255 50.475 0.715 ;
        RECT 50.645 0.085 50.915 0.545 ;
        RECT 51.085 0.255 51.415 0.715 ;
        RECT 51.585 0.085 51.835 0.885 ;
        RECT 0.000 -0.085 51.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 5.355 0.315 5.525 ;
        RECT 0.605 5.355 0.775 5.525 ;
        RECT 1.065 5.355 1.235 5.525 ;
        RECT 1.525 5.355 1.695 5.525 ;
        RECT 1.985 5.355 2.155 5.525 ;
        RECT 2.445 5.355 2.615 5.525 ;
        RECT 2.905 5.355 3.075 5.525 ;
        RECT 3.365 5.355 3.535 5.525 ;
        RECT 3.825 5.355 3.995 5.525 ;
        RECT 4.285 5.355 4.455 5.525 ;
        RECT 4.745 5.355 4.915 5.525 ;
        RECT 5.205 5.355 5.375 5.525 ;
        RECT 5.665 5.355 5.835 5.525 ;
        RECT 6.125 5.355 6.295 5.525 ;
        RECT 6.585 5.355 6.755 5.525 ;
        RECT 7.045 5.355 7.215 5.525 ;
        RECT 7.505 5.355 7.675 5.525 ;
        RECT 7.965 5.355 8.135 5.525 ;
        RECT 8.425 5.355 8.595 5.525 ;
        RECT 8.885 5.355 9.055 5.525 ;
        RECT 9.345 5.355 9.515 5.525 ;
        RECT 9.805 5.355 9.975 5.525 ;
        RECT 10.265 5.355 10.435 5.525 ;
        RECT 10.725 5.355 10.895 5.525 ;
        RECT 11.185 5.355 11.355 5.525 ;
        RECT 11.645 5.355 11.815 5.525 ;
        RECT 12.105 5.355 12.275 5.525 ;
        RECT 12.565 5.355 12.735 5.525 ;
        RECT 13.025 5.355 13.195 5.525 ;
        RECT 13.485 5.355 13.655 5.525 ;
        RECT 13.945 5.355 14.115 5.525 ;
        RECT 14.405 5.355 14.575 5.525 ;
        RECT 14.865 5.355 15.035 5.525 ;
        RECT 15.325 5.355 15.495 5.525 ;
        RECT 15.785 5.355 15.955 5.525 ;
        RECT 16.245 5.355 16.415 5.525 ;
        RECT 16.705 5.355 16.875 5.525 ;
        RECT 17.165 5.355 17.335 5.525 ;
        RECT 17.625 5.355 17.795 5.525 ;
        RECT 18.085 5.355 18.255 5.525 ;
        RECT 18.545 5.355 18.715 5.525 ;
        RECT 19.005 5.355 19.175 5.525 ;
        RECT 19.465 5.355 19.635 5.525 ;
        RECT 19.925 5.355 20.095 5.525 ;
        RECT 20.385 5.355 20.555 5.525 ;
        RECT 20.845 5.355 21.015 5.525 ;
        RECT 21.305 5.355 21.475 5.525 ;
        RECT 21.765 5.355 21.935 5.525 ;
        RECT 22.225 5.355 22.395 5.525 ;
        RECT 22.685 5.355 22.855 5.525 ;
        RECT 23.145 5.355 23.315 5.525 ;
        RECT 23.605 5.355 23.775 5.525 ;
        RECT 24.065 5.355 24.235 5.525 ;
        RECT 24.525 5.355 24.695 5.525 ;
        RECT 24.985 5.355 25.155 5.525 ;
        RECT 25.445 5.355 25.615 5.525 ;
        RECT 25.905 5.355 26.075 5.525 ;
        RECT 26.365 5.355 26.535 5.525 ;
        RECT 26.825 5.355 26.995 5.525 ;
        RECT 27.285 5.355 27.455 5.525 ;
        RECT 27.745 5.355 27.915 5.525 ;
        RECT 28.205 5.355 28.375 5.525 ;
        RECT 28.665 5.355 28.835 5.525 ;
        RECT 29.125 5.355 29.295 5.525 ;
        RECT 29.585 5.355 29.755 5.525 ;
        RECT 30.045 5.355 30.215 5.525 ;
        RECT 30.505 5.355 30.675 5.525 ;
        RECT 30.965 5.355 31.135 5.525 ;
        RECT 31.425 5.355 31.595 5.525 ;
        RECT 31.885 5.355 32.055 5.525 ;
        RECT 32.345 5.355 32.515 5.525 ;
        RECT 32.805 5.355 32.975 5.525 ;
        RECT 33.265 5.355 33.435 5.525 ;
        RECT 33.725 5.355 33.895 5.525 ;
        RECT 34.185 5.355 34.355 5.525 ;
        RECT 34.645 5.355 34.815 5.525 ;
        RECT 35.105 5.355 35.275 5.525 ;
        RECT 35.565 5.355 35.735 5.525 ;
        RECT 36.025 5.355 36.195 5.525 ;
        RECT 36.485 5.355 36.655 5.525 ;
        RECT 36.945 5.355 37.115 5.525 ;
        RECT 37.405 5.355 37.575 5.525 ;
        RECT 37.865 5.355 38.035 5.525 ;
        RECT 38.325 5.355 38.495 5.525 ;
        RECT 38.785 5.355 38.955 5.525 ;
        RECT 39.245 5.355 39.415 5.525 ;
        RECT 39.705 5.355 39.875 5.525 ;
        RECT 40.165 5.355 40.335 5.525 ;
        RECT 40.625 5.355 40.795 5.525 ;
        RECT 41.085 5.355 41.255 5.525 ;
        RECT 41.545 5.355 41.715 5.525 ;
        RECT 42.005 5.355 42.175 5.525 ;
        RECT 42.465 5.355 42.635 5.525 ;
        RECT 42.925 5.355 43.095 5.525 ;
        RECT 43.385 5.355 43.555 5.525 ;
        RECT 43.845 5.355 44.015 5.525 ;
        RECT 44.305 5.355 44.475 5.525 ;
        RECT 44.765 5.355 44.935 5.525 ;
        RECT 45.225 5.355 45.395 5.525 ;
        RECT 45.685 5.355 45.855 5.525 ;
        RECT 46.145 5.355 46.315 5.525 ;
        RECT 46.605 5.355 46.775 5.525 ;
        RECT 47.065 5.355 47.235 5.525 ;
        RECT 47.525 5.355 47.695 5.525 ;
        RECT 47.985 5.355 48.155 5.525 ;
        RECT 48.445 5.355 48.615 5.525 ;
        RECT 48.905 5.355 49.075 5.525 ;
        RECT 49.365 5.355 49.535 5.525 ;
        RECT 49.825 5.355 49.995 5.525 ;
        RECT 50.285 5.355 50.455 5.525 ;
        RECT 50.745 5.355 50.915 5.525 ;
        RECT 51.205 5.355 51.375 5.525 ;
        RECT 51.665 5.355 51.835 5.525 ;
        RECT 0.645 3.130 0.815 3.300 ;
        RECT 1.585 3.130 1.755 3.300 ;
        RECT 2.565 3.130 2.735 3.300 ;
        RECT 3.045 3.485 3.215 3.655 ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.645 2.140 0.815 2.310 ;
        RECT 1.585 2.140 1.755 2.310 ;
        RECT 2.565 2.140 2.735 2.310 ;
        RECT 3.515 3.130 3.685 3.300 ;
        RECT 3.985 3.485 4.155 3.655 ;
        RECT 3.045 1.785 3.215 1.955 ;
        RECT 3.515 2.140 3.685 2.310 ;
        RECT 4.465 3.130 4.635 3.300 ;
        RECT 8.245 3.130 8.415 3.300 ;
        RECT 8.725 3.485 8.895 3.655 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 3.985 1.785 4.155 1.955 ;
        RECT 4.465 2.140 4.635 2.310 ;
        RECT 8.245 2.140 8.415 2.310 ;
        RECT 9.195 3.130 9.365 3.300 ;
        RECT 9.665 3.485 9.835 3.655 ;
        RECT 8.725 1.785 8.895 1.955 ;
        RECT 9.195 2.140 9.365 2.310 ;
        RECT 10.145 3.130 10.315 3.300 ;
        RECT 11.125 3.130 11.295 3.300 ;
        RECT 12.065 3.130 12.235 3.300 ;
        RECT 13.525 3.130 13.695 3.300 ;
        RECT 14.465 3.130 14.635 3.300 ;
        RECT 15.445 3.130 15.615 3.300 ;
        RECT 15.925 3.485 16.095 3.655 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 14.405 2.635 14.575 2.805 ;
        RECT 14.865 2.635 15.035 2.805 ;
        RECT 15.325 2.635 15.495 2.805 ;
        RECT 9.665 1.785 9.835 1.955 ;
        RECT 10.145 2.140 10.315 2.310 ;
        RECT 11.125 2.140 11.295 2.310 ;
        RECT 12.065 2.140 12.235 2.310 ;
        RECT 13.525 2.140 13.695 2.310 ;
        RECT 14.465 2.140 14.635 2.310 ;
        RECT 15.445 2.140 15.615 2.310 ;
        RECT 16.395 3.130 16.565 3.300 ;
        RECT 16.865 3.485 17.035 3.655 ;
        RECT 15.925 1.785 16.095 1.955 ;
        RECT 16.395 2.140 16.565 2.310 ;
        RECT 17.345 3.130 17.515 3.300 ;
        RECT 21.125 3.130 21.295 3.300 ;
        RECT 21.605 3.485 21.775 3.655 ;
        RECT 17.625 2.635 17.795 2.805 ;
        RECT 18.085 2.635 18.255 2.805 ;
        RECT 18.545 2.635 18.715 2.805 ;
        RECT 19.005 2.635 19.175 2.805 ;
        RECT 19.465 2.635 19.635 2.805 ;
        RECT 19.925 2.635 20.095 2.805 ;
        RECT 20.385 2.635 20.555 2.805 ;
        RECT 20.845 2.635 21.015 2.805 ;
        RECT 16.865 1.785 17.035 1.955 ;
        RECT 17.345 2.140 17.515 2.310 ;
        RECT 21.125 2.140 21.295 2.310 ;
        RECT 22.075 3.130 22.245 3.300 ;
        RECT 22.545 3.485 22.715 3.655 ;
        RECT 21.605 1.785 21.775 1.955 ;
        RECT 22.075 2.140 22.245 2.310 ;
        RECT 23.025 3.130 23.195 3.300 ;
        RECT 24.005 3.130 24.175 3.300 ;
        RECT 24.945 3.130 25.115 3.300 ;
        RECT 26.865 3.130 27.035 3.300 ;
        RECT 27.805 3.130 27.975 3.300 ;
        RECT 28.785 3.130 28.955 3.300 ;
        RECT 29.265 3.485 29.435 3.655 ;
        RECT 23.145 2.635 23.315 2.805 ;
        RECT 23.605 2.635 23.775 2.805 ;
        RECT 24.065 2.635 24.235 2.805 ;
        RECT 24.525 2.635 24.695 2.805 ;
        RECT 24.985 2.635 25.155 2.805 ;
        RECT 25.445 2.635 25.615 2.805 ;
        RECT 25.905 2.635 26.075 2.805 ;
        RECT 26.365 2.635 26.535 2.805 ;
        RECT 26.825 2.635 26.995 2.805 ;
        RECT 27.285 2.635 27.455 2.805 ;
        RECT 27.745 2.635 27.915 2.805 ;
        RECT 28.205 2.635 28.375 2.805 ;
        RECT 28.665 2.635 28.835 2.805 ;
        RECT 22.545 1.785 22.715 1.955 ;
        RECT 23.025 2.140 23.195 2.310 ;
        RECT 24.005 2.140 24.175 2.310 ;
        RECT 24.945 2.140 25.115 2.310 ;
        RECT 26.865 2.140 27.035 2.310 ;
        RECT 27.805 2.140 27.975 2.310 ;
        RECT 28.785 2.140 28.955 2.310 ;
        RECT 29.735 3.130 29.905 3.300 ;
        RECT 30.205 3.485 30.375 3.655 ;
        RECT 29.265 1.785 29.435 1.955 ;
        RECT 29.735 2.140 29.905 2.310 ;
        RECT 30.685 3.130 30.855 3.300 ;
        RECT 34.465 3.130 34.635 3.300 ;
        RECT 34.945 3.485 35.115 3.655 ;
        RECT 30.965 2.635 31.135 2.805 ;
        RECT 31.425 2.635 31.595 2.805 ;
        RECT 31.885 2.635 32.055 2.805 ;
        RECT 32.345 2.635 32.515 2.805 ;
        RECT 32.805 2.635 32.975 2.805 ;
        RECT 33.265 2.635 33.435 2.805 ;
        RECT 33.725 2.635 33.895 2.805 ;
        RECT 34.185 2.635 34.355 2.805 ;
        RECT 30.205 1.785 30.375 1.955 ;
        RECT 30.685 2.140 30.855 2.310 ;
        RECT 34.465 2.140 34.635 2.310 ;
        RECT 35.415 3.130 35.585 3.300 ;
        RECT 35.885 3.485 36.055 3.655 ;
        RECT 34.945 1.785 35.115 1.955 ;
        RECT 35.415 2.140 35.585 2.310 ;
        RECT 36.365 3.130 36.535 3.300 ;
        RECT 37.345 3.130 37.515 3.300 ;
        RECT 38.285 3.130 38.455 3.300 ;
        RECT 39.745 3.130 39.915 3.300 ;
        RECT 40.685 3.130 40.855 3.300 ;
        RECT 41.665 3.130 41.835 3.300 ;
        RECT 42.145 3.485 42.315 3.655 ;
        RECT 36.485 2.635 36.655 2.805 ;
        RECT 36.945 2.635 37.115 2.805 ;
        RECT 37.405 2.635 37.575 2.805 ;
        RECT 37.865 2.635 38.035 2.805 ;
        RECT 38.325 2.635 38.495 2.805 ;
        RECT 38.785 2.635 38.955 2.805 ;
        RECT 39.245 2.635 39.415 2.805 ;
        RECT 39.705 2.635 39.875 2.805 ;
        RECT 40.165 2.635 40.335 2.805 ;
        RECT 40.625 2.635 40.795 2.805 ;
        RECT 41.085 2.635 41.255 2.805 ;
        RECT 41.545 2.635 41.715 2.805 ;
        RECT 35.885 1.785 36.055 1.955 ;
        RECT 36.365 2.140 36.535 2.310 ;
        RECT 37.345 2.140 37.515 2.310 ;
        RECT 38.285 2.140 38.455 2.310 ;
        RECT 39.745 2.140 39.915 2.310 ;
        RECT 40.685 2.140 40.855 2.310 ;
        RECT 41.665 2.140 41.835 2.310 ;
        RECT 42.615 3.130 42.785 3.300 ;
        RECT 43.085 3.485 43.255 3.655 ;
        RECT 42.145 1.785 42.315 1.955 ;
        RECT 42.615 2.140 42.785 2.310 ;
        RECT 43.565 3.130 43.735 3.300 ;
        RECT 47.345 3.130 47.515 3.300 ;
        RECT 47.825 3.485 47.995 3.655 ;
        RECT 43.845 2.635 44.015 2.805 ;
        RECT 44.305 2.635 44.475 2.805 ;
        RECT 44.765 2.635 44.935 2.805 ;
        RECT 45.225 2.635 45.395 2.805 ;
        RECT 45.685 2.635 45.855 2.805 ;
        RECT 46.145 2.635 46.315 2.805 ;
        RECT 46.605 2.635 46.775 2.805 ;
        RECT 47.065 2.635 47.235 2.805 ;
        RECT 43.085 1.785 43.255 1.955 ;
        RECT 43.565 2.140 43.735 2.310 ;
        RECT 47.345 2.140 47.515 2.310 ;
        RECT 48.295 3.130 48.465 3.300 ;
        RECT 48.765 3.485 48.935 3.655 ;
        RECT 47.825 1.785 47.995 1.955 ;
        RECT 48.295 2.140 48.465 2.310 ;
        RECT 49.245 3.130 49.415 3.300 ;
        RECT 50.225 3.130 50.395 3.300 ;
        RECT 51.165 3.130 51.335 3.300 ;
        RECT 49.365 2.635 49.535 2.805 ;
        RECT 49.825 2.635 49.995 2.805 ;
        RECT 50.285 2.635 50.455 2.805 ;
        RECT 50.745 2.635 50.915 2.805 ;
        RECT 51.205 2.635 51.375 2.805 ;
        RECT 51.665 2.635 51.835 2.805 ;
        RECT 48.765 1.785 48.935 1.955 ;
        RECT 49.245 2.140 49.415 2.310 ;
        RECT 50.225 2.140 50.395 2.310 ;
        RECT 51.165 2.140 51.335 2.310 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
        RECT 14.405 -0.085 14.575 0.085 ;
        RECT 14.865 -0.085 15.035 0.085 ;
        RECT 15.325 -0.085 15.495 0.085 ;
        RECT 15.785 -0.085 15.955 0.085 ;
        RECT 16.245 -0.085 16.415 0.085 ;
        RECT 16.705 -0.085 16.875 0.085 ;
        RECT 17.165 -0.085 17.335 0.085 ;
        RECT 17.625 -0.085 17.795 0.085 ;
        RECT 18.085 -0.085 18.255 0.085 ;
        RECT 18.545 -0.085 18.715 0.085 ;
        RECT 19.005 -0.085 19.175 0.085 ;
        RECT 19.465 -0.085 19.635 0.085 ;
        RECT 19.925 -0.085 20.095 0.085 ;
        RECT 20.385 -0.085 20.555 0.085 ;
        RECT 20.845 -0.085 21.015 0.085 ;
        RECT 21.305 -0.085 21.475 0.085 ;
        RECT 21.765 -0.085 21.935 0.085 ;
        RECT 22.225 -0.085 22.395 0.085 ;
        RECT 22.685 -0.085 22.855 0.085 ;
        RECT 23.145 -0.085 23.315 0.085 ;
        RECT 23.605 -0.085 23.775 0.085 ;
        RECT 24.065 -0.085 24.235 0.085 ;
        RECT 24.525 -0.085 24.695 0.085 ;
        RECT 24.985 -0.085 25.155 0.085 ;
        RECT 25.445 -0.085 25.615 0.085 ;
        RECT 25.905 -0.085 26.075 0.085 ;
        RECT 26.365 -0.085 26.535 0.085 ;
        RECT 26.825 -0.085 26.995 0.085 ;
        RECT 27.285 -0.085 27.455 0.085 ;
        RECT 27.745 -0.085 27.915 0.085 ;
        RECT 28.205 -0.085 28.375 0.085 ;
        RECT 28.665 -0.085 28.835 0.085 ;
        RECT 29.125 -0.085 29.295 0.085 ;
        RECT 29.585 -0.085 29.755 0.085 ;
        RECT 30.045 -0.085 30.215 0.085 ;
        RECT 30.505 -0.085 30.675 0.085 ;
        RECT 30.965 -0.085 31.135 0.085 ;
        RECT 31.425 -0.085 31.595 0.085 ;
        RECT 31.885 -0.085 32.055 0.085 ;
        RECT 32.345 -0.085 32.515 0.085 ;
        RECT 32.805 -0.085 32.975 0.085 ;
        RECT 33.265 -0.085 33.435 0.085 ;
        RECT 33.725 -0.085 33.895 0.085 ;
        RECT 34.185 -0.085 34.355 0.085 ;
        RECT 34.645 -0.085 34.815 0.085 ;
        RECT 35.105 -0.085 35.275 0.085 ;
        RECT 35.565 -0.085 35.735 0.085 ;
        RECT 36.025 -0.085 36.195 0.085 ;
        RECT 36.485 -0.085 36.655 0.085 ;
        RECT 36.945 -0.085 37.115 0.085 ;
        RECT 37.405 -0.085 37.575 0.085 ;
        RECT 37.865 -0.085 38.035 0.085 ;
        RECT 38.325 -0.085 38.495 0.085 ;
        RECT 38.785 -0.085 38.955 0.085 ;
        RECT 39.245 -0.085 39.415 0.085 ;
        RECT 39.705 -0.085 39.875 0.085 ;
        RECT 40.165 -0.085 40.335 0.085 ;
        RECT 40.625 -0.085 40.795 0.085 ;
        RECT 41.085 -0.085 41.255 0.085 ;
        RECT 41.545 -0.085 41.715 0.085 ;
        RECT 42.005 -0.085 42.175 0.085 ;
        RECT 42.465 -0.085 42.635 0.085 ;
        RECT 42.925 -0.085 43.095 0.085 ;
        RECT 43.385 -0.085 43.555 0.085 ;
        RECT 43.845 -0.085 44.015 0.085 ;
        RECT 44.305 -0.085 44.475 0.085 ;
        RECT 44.765 -0.085 44.935 0.085 ;
        RECT 45.225 -0.085 45.395 0.085 ;
        RECT 45.685 -0.085 45.855 0.085 ;
        RECT 46.145 -0.085 46.315 0.085 ;
        RECT 46.605 -0.085 46.775 0.085 ;
        RECT 47.065 -0.085 47.235 0.085 ;
        RECT 47.525 -0.085 47.695 0.085 ;
        RECT 47.985 -0.085 48.155 0.085 ;
        RECT 48.445 -0.085 48.615 0.085 ;
        RECT 48.905 -0.085 49.075 0.085 ;
        RECT 49.365 -0.085 49.535 0.085 ;
        RECT 49.825 -0.085 49.995 0.085 ;
        RECT 50.285 -0.085 50.455 0.085 ;
        RECT 50.745 -0.085 50.915 0.085 ;
        RECT 51.205 -0.085 51.375 0.085 ;
        RECT 51.665 -0.085 51.835 0.085 ;
      LAYER met1 ;
        RECT 0.585 3.285 0.875 3.330 ;
        RECT 1.525 3.285 1.815 3.330 ;
        RECT 2.505 3.285 2.795 3.330 ;
        RECT 3.455 3.285 3.745 3.330 ;
        RECT 4.405 3.285 4.695 3.330 ;
        RECT 0.585 3.145 4.695 3.285 ;
        RECT 0.585 3.100 0.875 3.145 ;
        RECT 1.525 3.100 1.815 3.145 ;
        RECT 2.505 3.100 2.795 3.145 ;
        RECT 3.455 3.100 3.745 3.145 ;
        RECT 4.405 3.100 4.695 3.145 ;
        RECT 8.185 3.285 8.475 3.330 ;
        RECT 9.135 3.285 9.425 3.330 ;
        RECT 10.085 3.285 10.375 3.330 ;
        RECT 11.065 3.285 11.355 3.330 ;
        RECT 12.005 3.285 12.295 3.330 ;
        RECT 8.185 3.145 12.295 3.285 ;
        RECT 8.185 3.100 8.475 3.145 ;
        RECT 9.135 3.100 9.425 3.145 ;
        RECT 10.085 3.100 10.375 3.145 ;
        RECT 11.065 3.100 11.355 3.145 ;
        RECT 12.005 3.100 12.295 3.145 ;
        RECT 13.465 3.285 13.755 3.330 ;
        RECT 14.405 3.285 14.695 3.330 ;
        RECT 15.385 3.285 15.675 3.330 ;
        RECT 16.335 3.285 16.625 3.330 ;
        RECT 17.285 3.285 17.575 3.330 ;
        RECT 13.465 3.145 17.575 3.285 ;
        RECT 13.465 3.100 13.755 3.145 ;
        RECT 14.405 3.100 14.695 3.145 ;
        RECT 15.385 3.100 15.675 3.145 ;
        RECT 16.335 3.100 16.625 3.145 ;
        RECT 17.285 3.100 17.575 3.145 ;
        RECT 21.065 3.285 21.355 3.330 ;
        RECT 22.015 3.285 22.305 3.330 ;
        RECT 22.965 3.285 23.255 3.330 ;
        RECT 23.945 3.285 24.235 3.330 ;
        RECT 24.885 3.285 25.175 3.330 ;
        RECT 21.065 3.145 25.175 3.285 ;
        RECT 21.065 3.100 21.355 3.145 ;
        RECT 22.015 3.100 22.305 3.145 ;
        RECT 22.965 3.100 23.255 3.145 ;
        RECT 23.945 3.100 24.235 3.145 ;
        RECT 24.885 3.100 25.175 3.145 ;
        RECT 26.805 3.285 27.095 3.330 ;
        RECT 27.745 3.285 28.035 3.330 ;
        RECT 28.725 3.285 29.015 3.330 ;
        RECT 29.675 3.285 29.965 3.330 ;
        RECT 30.625 3.285 30.915 3.330 ;
        RECT 26.805 3.145 30.915 3.285 ;
        RECT 26.805 3.100 27.095 3.145 ;
        RECT 27.745 3.100 28.035 3.145 ;
        RECT 28.725 3.100 29.015 3.145 ;
        RECT 29.675 3.100 29.965 3.145 ;
        RECT 30.625 3.100 30.915 3.145 ;
        RECT 34.405 3.285 34.695 3.330 ;
        RECT 35.355 3.285 35.645 3.330 ;
        RECT 36.305 3.285 36.595 3.330 ;
        RECT 37.285 3.285 37.575 3.330 ;
        RECT 38.225 3.285 38.515 3.330 ;
        RECT 34.405 3.145 38.515 3.285 ;
        RECT 34.405 3.100 34.695 3.145 ;
        RECT 35.355 3.100 35.645 3.145 ;
        RECT 36.305 3.100 36.595 3.145 ;
        RECT 37.285 3.100 37.575 3.145 ;
        RECT 38.225 3.100 38.515 3.145 ;
        RECT 39.685 3.285 39.975 3.330 ;
        RECT 40.625 3.285 40.915 3.330 ;
        RECT 41.605 3.285 41.895 3.330 ;
        RECT 42.555 3.285 42.845 3.330 ;
        RECT 43.505 3.285 43.795 3.330 ;
        RECT 39.685 3.145 43.795 3.285 ;
        RECT 39.685 3.100 39.975 3.145 ;
        RECT 40.625 3.100 40.915 3.145 ;
        RECT 41.605 3.100 41.895 3.145 ;
        RECT 42.555 3.100 42.845 3.145 ;
        RECT 43.505 3.100 43.795 3.145 ;
        RECT 47.285 3.285 47.575 3.330 ;
        RECT 48.235 3.285 48.525 3.330 ;
        RECT 49.185 3.285 49.475 3.330 ;
        RECT 50.165 3.285 50.455 3.330 ;
        RECT 51.105 3.285 51.395 3.330 ;
        RECT 47.285 3.145 51.395 3.285 ;
        RECT 47.285 3.100 47.575 3.145 ;
        RECT 48.235 3.100 48.525 3.145 ;
        RECT 49.185 3.100 49.475 3.145 ;
        RECT 50.165 3.100 50.455 3.145 ;
        RECT 51.105 3.100 51.395 3.145 ;
        RECT 0.585 2.295 0.875 2.340 ;
        RECT 1.525 2.295 1.815 2.340 ;
        RECT 2.505 2.295 2.795 2.340 ;
        RECT 3.455 2.295 3.745 2.340 ;
        RECT 4.405 2.295 4.695 2.340 ;
        RECT 0.585 2.155 4.695 2.295 ;
        RECT 0.585 2.110 0.875 2.155 ;
        RECT 1.525 2.110 1.815 2.155 ;
        RECT 2.505 2.110 2.795 2.155 ;
        RECT 3.455 2.110 3.745 2.155 ;
        RECT 4.405 2.110 4.695 2.155 ;
        RECT 8.185 2.295 8.475 2.340 ;
        RECT 9.135 2.295 9.425 2.340 ;
        RECT 10.085 2.295 10.375 2.340 ;
        RECT 11.065 2.295 11.355 2.340 ;
        RECT 12.005 2.295 12.295 2.340 ;
        RECT 8.185 2.155 12.295 2.295 ;
        RECT 8.185 2.110 8.475 2.155 ;
        RECT 9.135 2.110 9.425 2.155 ;
        RECT 10.085 2.110 10.375 2.155 ;
        RECT 11.065 2.110 11.355 2.155 ;
        RECT 12.005 2.110 12.295 2.155 ;
        RECT 13.465 2.295 13.755 2.340 ;
        RECT 14.405 2.295 14.695 2.340 ;
        RECT 15.385 2.295 15.675 2.340 ;
        RECT 16.335 2.295 16.625 2.340 ;
        RECT 17.285 2.295 17.575 2.340 ;
        RECT 13.465 2.155 17.575 2.295 ;
        RECT 13.465 2.110 13.755 2.155 ;
        RECT 14.405 2.110 14.695 2.155 ;
        RECT 15.385 2.110 15.675 2.155 ;
        RECT 16.335 2.110 16.625 2.155 ;
        RECT 17.285 2.110 17.575 2.155 ;
        RECT 21.065 2.295 21.355 2.340 ;
        RECT 22.015 2.295 22.305 2.340 ;
        RECT 22.965 2.295 23.255 2.340 ;
        RECT 23.945 2.295 24.235 2.340 ;
        RECT 24.885 2.295 25.175 2.340 ;
        RECT 21.065 2.155 25.175 2.295 ;
        RECT 21.065 2.110 21.355 2.155 ;
        RECT 22.015 2.110 22.305 2.155 ;
        RECT 22.965 2.110 23.255 2.155 ;
        RECT 23.945 2.110 24.235 2.155 ;
        RECT 24.885 2.110 25.175 2.155 ;
        RECT 26.805 2.295 27.095 2.340 ;
        RECT 27.745 2.295 28.035 2.340 ;
        RECT 28.725 2.295 29.015 2.340 ;
        RECT 29.675 2.295 29.965 2.340 ;
        RECT 30.625 2.295 30.915 2.340 ;
        RECT 26.805 2.155 30.915 2.295 ;
        RECT 26.805 2.110 27.095 2.155 ;
        RECT 27.745 2.110 28.035 2.155 ;
        RECT 28.725 2.110 29.015 2.155 ;
        RECT 29.675 2.110 29.965 2.155 ;
        RECT 30.625 2.110 30.915 2.155 ;
        RECT 34.405 2.295 34.695 2.340 ;
        RECT 35.355 2.295 35.645 2.340 ;
        RECT 36.305 2.295 36.595 2.340 ;
        RECT 37.285 2.295 37.575 2.340 ;
        RECT 38.225 2.295 38.515 2.340 ;
        RECT 34.405 2.155 38.515 2.295 ;
        RECT 34.405 2.110 34.695 2.155 ;
        RECT 35.355 2.110 35.645 2.155 ;
        RECT 36.305 2.110 36.595 2.155 ;
        RECT 37.285 2.110 37.575 2.155 ;
        RECT 38.225 2.110 38.515 2.155 ;
        RECT 39.685 2.295 39.975 2.340 ;
        RECT 40.625 2.295 40.915 2.340 ;
        RECT 41.605 2.295 41.895 2.340 ;
        RECT 42.555 2.295 42.845 2.340 ;
        RECT 43.505 2.295 43.795 2.340 ;
        RECT 39.685 2.155 43.795 2.295 ;
        RECT 39.685 2.110 39.975 2.155 ;
        RECT 40.625 2.110 40.915 2.155 ;
        RECT 41.605 2.110 41.895 2.155 ;
        RECT 42.555 2.110 42.845 2.155 ;
        RECT 43.505 2.110 43.795 2.155 ;
        RECT 47.285 2.295 47.575 2.340 ;
        RECT 48.235 2.295 48.525 2.340 ;
        RECT 49.185 2.295 49.475 2.340 ;
        RECT 50.165 2.295 50.455 2.340 ;
        RECT 51.105 2.295 51.395 2.340 ;
        RECT 47.285 2.155 51.395 2.295 ;
        RECT 47.285 2.110 47.575 2.155 ;
        RECT 48.235 2.110 48.525 2.155 ;
        RECT 49.185 2.110 49.475 2.155 ;
        RECT 50.165 2.110 50.455 2.155 ;
        RECT 51.105 2.110 51.395 2.155 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__muxb16to1_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__nand2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.990 1.075 1.375 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.055 0.430 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.025 0.105 1.475 1.015 ;
        RECT 0.140 -0.085 0.310 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.491500 ;
    PORT
      LAYER li1 ;
        RECT 0.535 1.485 0.915 2.465 ;
        RECT 0.650 0.885 0.820 1.485 ;
        RECT 0.650 0.255 1.395 0.885 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.840 2.805 ;
        RECT 0.085 1.495 0.365 2.635 ;
        RECT 1.135 1.495 1.395 2.635 ;
        RECT 0.085 0.085 0.395 0.885 ;
        RECT 0.000 -0.085 1.840 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand2_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__nand2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.075 1.780 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.895 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.395 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.820500 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.665 0.895 2.465 ;
        RECT 1.455 1.665 1.835 2.465 ;
        RECT 0.515 1.495 2.230 1.665 ;
        RECT 1.950 0.905 2.230 1.495 ;
        RECT 1.455 0.655 2.230 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.085 1.495 0.345 2.635 ;
        RECT 1.115 1.835 1.285 2.635 ;
        RECT 2.055 1.835 2.310 2.635 ;
        RECT 0.085 0.715 1.285 0.885 ;
        RECT 0.085 0.255 0.425 0.715 ;
        RECT 0.645 0.085 0.815 0.545 ;
        RECT 0.985 0.485 1.285 0.715 ;
        RECT 0.985 0.255 2.305 0.485 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand2_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__nand2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 2.865 1.075 4.115 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.110 1.075 1.880 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.275 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.608500 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.665 0.895 2.465 ;
        RECT 1.455 1.665 1.835 2.465 ;
        RECT 2.395 1.665 2.775 2.465 ;
        RECT 3.335 1.665 3.715 2.465 ;
        RECT 0.515 1.495 3.715 1.665 ;
        RECT 2.395 0.805 2.695 1.495 ;
        RECT 2.395 0.635 3.715 0.805 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.090 1.495 0.345 2.635 ;
        RECT 1.115 1.835 1.285 2.635 ;
        RECT 2.055 1.835 2.225 2.635 ;
        RECT 2.995 1.835 3.165 2.635 ;
        RECT 3.935 1.835 4.185 2.635 ;
        RECT 0.090 0.715 2.225 0.905 ;
        RECT 0.090 0.255 0.425 0.715 ;
        RECT 0.645 0.085 0.815 0.545 ;
        RECT 0.985 0.255 1.365 0.715 ;
        RECT 1.585 0.085 1.755 0.545 ;
        RECT 1.925 0.465 2.225 0.715 ;
        RECT 3.935 0.465 4.185 0.885 ;
        RECT 1.925 0.255 4.185 0.465 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand2_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__nand2_6
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand2_6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.665000 ;
    PORT
      LAYER li1 ;
        RECT 3.805 1.055 5.155 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.665000 ;
    PORT
      LAYER li1 ;
        RECT 0.395 1.055 2.765 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 6.155 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.429000 ;
    PORT
      LAYER li1 ;
        RECT 0.565 1.665 0.895 2.465 ;
        RECT 1.505 1.665 1.835 2.465 ;
        RECT 2.445 1.665 2.775 2.465 ;
        RECT 3.385 1.665 3.715 2.465 ;
        RECT 4.325 1.665 4.655 2.465 ;
        RECT 5.265 1.665 5.595 2.465 ;
        RECT 0.565 1.495 5.595 1.665 ;
        RECT 3.335 0.885 3.635 1.495 ;
        RECT 5.325 1.325 5.595 1.495 ;
        RECT 5.325 1.055 5.915 1.325 ;
        RECT 5.325 0.885 5.595 1.055 ;
        RECT 3.335 0.635 5.595 0.885 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.125 1.495 0.395 2.635 ;
        RECT 1.065 1.835 1.335 2.635 ;
        RECT 2.005 1.835 2.275 2.635 ;
        RECT 2.945 1.835 3.215 2.635 ;
        RECT 3.885 1.835 4.155 2.635 ;
        RECT 4.825 1.835 5.095 2.635 ;
        RECT 5.765 1.495 6.035 2.635 ;
        RECT 0.090 0.715 3.165 0.885 ;
        RECT 0.090 0.255 0.425 0.715 ;
        RECT 0.595 0.085 0.865 0.545 ;
        RECT 1.035 0.255 1.365 0.715 ;
        RECT 1.535 0.085 1.805 0.545 ;
        RECT 1.975 0.255 2.305 0.715 ;
        RECT 2.475 0.085 2.745 0.545 ;
        RECT 2.915 0.465 3.165 0.715 ;
        RECT 5.765 0.465 6.065 0.885 ;
        RECT 2.915 0.255 6.065 0.465 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand2_6

#--------EOF---------

MACRO sky130_fd_sc_hdll__nand2_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand2_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.280 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.220000 ;
    PORT
      LAYER li1 ;
        RECT 4.740 1.075 7.005 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.220000 ;
    PORT
      LAYER li1 ;
        RECT 0.510 1.075 3.715 1.295 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.280 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 8.155 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.470 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.280 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.184500 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.665 0.895 2.465 ;
        RECT 1.455 1.665 1.835 2.465 ;
        RECT 2.395 1.665 2.775 2.465 ;
        RECT 3.335 1.665 3.715 2.465 ;
        RECT 4.275 1.665 4.655 2.465 ;
        RECT 5.215 1.665 5.595 2.465 ;
        RECT 6.155 1.665 6.535 2.465 ;
        RECT 7.095 1.665 7.475 2.465 ;
        RECT 0.515 1.465 7.475 1.665 ;
        RECT 4.040 1.075 4.570 1.465 ;
        RECT 4.275 0.905 4.570 1.075 ;
        RECT 7.225 0.905 7.475 1.465 ;
        RECT 4.275 0.655 7.475 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.280 2.805 ;
        RECT 0.090 1.495 0.345 2.635 ;
        RECT 1.115 1.835 1.285 2.635 ;
        RECT 2.055 1.835 2.225 2.635 ;
        RECT 2.995 1.835 3.165 2.635 ;
        RECT 3.935 1.835 4.105 2.635 ;
        RECT 4.875 1.835 5.045 2.635 ;
        RECT 5.815 1.835 5.985 2.635 ;
        RECT 6.755 1.835 6.925 2.635 ;
        RECT 7.715 1.495 8.070 2.635 ;
        RECT 0.090 0.735 4.105 0.905 ;
        RECT 0.090 0.255 0.425 0.735 ;
        RECT 0.645 0.085 0.815 0.565 ;
        RECT 0.985 0.255 1.365 0.735 ;
        RECT 1.585 0.085 1.755 0.565 ;
        RECT 1.925 0.255 2.305 0.735 ;
        RECT 2.525 0.085 2.695 0.565 ;
        RECT 2.865 0.255 3.245 0.735 ;
        RECT 3.465 0.085 3.635 0.565 ;
        RECT 3.805 0.485 4.105 0.735 ;
        RECT 7.695 0.485 8.070 0.905 ;
        RECT 3.805 0.255 8.070 0.485 ;
        RECT 0.000 -0.085 8.280 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand2_8

#--------EOF---------

MACRO sky130_fd_sc_hdll__nand2_12
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand2_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.960 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.330000 ;
    PORT
      LAYER li1 ;
        RECT 6.625 1.055 10.695 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.330000 ;
    PORT
      LAYER li1 ;
        RECT 0.335 1.055 5.765 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.960 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 11.795 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 12.150 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.960 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.858000 ;
    PORT
      LAYER li1 ;
        RECT 0.565 1.665 0.895 2.465 ;
        RECT 1.505 1.665 1.835 2.465 ;
        RECT 2.445 1.665 2.775 2.465 ;
        RECT 3.385 1.665 3.715 2.465 ;
        RECT 4.325 1.665 4.655 2.465 ;
        RECT 5.265 1.665 5.595 2.465 ;
        RECT 6.205 1.665 6.535 2.465 ;
        RECT 7.145 1.665 7.475 2.465 ;
        RECT 8.085 1.665 8.415 2.465 ;
        RECT 9.025 1.665 9.355 2.465 ;
        RECT 9.965 1.665 10.295 2.465 ;
        RECT 10.905 1.665 11.235 2.465 ;
        RECT 0.565 1.495 11.235 1.665 ;
        RECT 6.045 1.055 6.455 1.495 ;
        RECT 6.155 0.885 6.455 1.055 ;
        RECT 10.965 1.325 11.235 1.495 ;
        RECT 10.965 1.055 11.435 1.325 ;
        RECT 10.965 0.885 11.235 1.055 ;
        RECT 6.155 0.635 11.235 0.885 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 11.960 2.805 ;
        RECT 0.125 1.495 0.395 2.635 ;
        RECT 1.065 1.835 1.335 2.635 ;
        RECT 2.005 1.835 2.275 2.635 ;
        RECT 2.945 1.835 3.215 2.635 ;
        RECT 3.885 1.835 4.155 2.635 ;
        RECT 4.825 1.835 5.095 2.635 ;
        RECT 5.765 1.835 6.035 2.635 ;
        RECT 6.705 1.835 6.975 2.635 ;
        RECT 7.645 1.835 7.915 2.635 ;
        RECT 8.585 1.835 8.855 2.635 ;
        RECT 9.525 1.835 9.795 2.635 ;
        RECT 10.465 1.835 10.735 2.635 ;
        RECT 11.405 1.495 11.675 2.635 ;
        RECT 0.090 0.715 5.985 0.885 ;
        RECT 0.090 0.255 0.425 0.715 ;
        RECT 0.595 0.085 0.865 0.545 ;
        RECT 1.035 0.255 1.365 0.715 ;
        RECT 1.535 0.085 1.805 0.545 ;
        RECT 1.975 0.255 2.305 0.715 ;
        RECT 2.475 0.085 2.745 0.545 ;
        RECT 2.915 0.255 3.245 0.715 ;
        RECT 3.415 0.085 3.685 0.545 ;
        RECT 3.855 0.255 4.185 0.715 ;
        RECT 4.355 0.085 4.625 0.545 ;
        RECT 4.795 0.255 5.125 0.715 ;
        RECT 5.295 0.085 5.565 0.545 ;
        RECT 5.735 0.465 5.985 0.715 ;
        RECT 11.455 0.465 11.705 0.885 ;
        RECT 5.735 0.255 11.705 0.465 ;
        RECT 0.000 -0.085 11.960 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand2_12

#--------EOF---------

MACRO sky130_fd_sc_hdll__nand2_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand2_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.640 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.440000 ;
    PORT
      LAYER li1 ;
        RECT 8.505 1.055 14.275 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.440000 ;
    PORT
      LAYER li1 ;
        RECT 0.395 1.055 7.525 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 15.640 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 15.555 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 15.830 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 15.640 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.499000 ;
    PORT
      LAYER li1 ;
        RECT 0.565 1.665 0.895 2.465 ;
        RECT 1.505 1.665 1.835 2.465 ;
        RECT 2.445 1.665 2.775 2.465 ;
        RECT 3.385 1.665 3.715 2.465 ;
        RECT 4.325 1.665 4.655 2.465 ;
        RECT 5.265 1.665 5.595 2.465 ;
        RECT 6.205 1.665 6.535 2.465 ;
        RECT 7.145 1.665 7.475 2.465 ;
        RECT 8.085 1.665 8.415 2.465 ;
        RECT 9.025 1.665 9.355 2.465 ;
        RECT 9.965 1.665 10.295 2.465 ;
        RECT 10.905 1.665 11.235 2.465 ;
        RECT 11.845 1.665 12.175 2.465 ;
        RECT 12.785 1.665 13.115 2.465 ;
        RECT 13.725 1.665 14.055 2.465 ;
        RECT 14.665 1.665 14.995 2.465 ;
        RECT 0.565 1.495 14.995 1.665 ;
        RECT 7.925 1.055 8.335 1.495 ;
        RECT 8.035 0.885 8.335 1.055 ;
        RECT 14.725 1.325 14.995 1.495 ;
        RECT 14.725 1.055 15.115 1.325 ;
        RECT 14.725 0.885 14.995 1.055 ;
        RECT 8.035 0.635 14.995 0.885 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 15.640 2.805 ;
        RECT 0.125 1.495 0.395 2.635 ;
        RECT 1.065 1.835 1.335 2.635 ;
        RECT 2.005 1.835 2.275 2.635 ;
        RECT 2.945 1.835 3.215 2.635 ;
        RECT 3.885 1.835 4.155 2.635 ;
        RECT 4.825 1.835 5.095 2.635 ;
        RECT 5.765 1.835 6.035 2.635 ;
        RECT 6.705 1.835 6.975 2.635 ;
        RECT 7.645 1.835 7.915 2.635 ;
        RECT 8.585 1.835 8.855 2.635 ;
        RECT 9.525 1.835 9.795 2.635 ;
        RECT 10.465 1.835 10.735 2.635 ;
        RECT 11.405 1.835 11.675 2.635 ;
        RECT 12.345 1.835 12.615 2.635 ;
        RECT 13.285 1.835 13.555 2.635 ;
        RECT 14.225 1.835 14.495 2.635 ;
        RECT 15.165 1.495 15.435 2.635 ;
        RECT 0.095 0.715 7.865 0.885 ;
        RECT 0.095 0.255 0.425 0.715 ;
        RECT 0.595 0.085 0.865 0.545 ;
        RECT 1.035 0.255 1.365 0.715 ;
        RECT 1.535 0.085 1.805 0.545 ;
        RECT 1.975 0.255 2.305 0.715 ;
        RECT 2.475 0.085 2.745 0.545 ;
        RECT 2.915 0.255 3.245 0.715 ;
        RECT 3.415 0.085 3.685 0.545 ;
        RECT 3.855 0.255 4.185 0.715 ;
        RECT 4.355 0.085 4.625 0.545 ;
        RECT 4.795 0.255 5.125 0.715 ;
        RECT 5.295 0.085 5.565 0.545 ;
        RECT 5.735 0.255 6.065 0.715 ;
        RECT 6.235 0.085 6.505 0.545 ;
        RECT 6.675 0.255 7.005 0.715 ;
        RECT 7.175 0.085 7.445 0.545 ;
        RECT 7.615 0.465 7.865 0.715 ;
        RECT 15.215 0.465 15.465 0.885 ;
        RECT 7.615 0.255 15.465 0.465 ;
        RECT 0.000 -0.085 15.640 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 14.405 2.635 14.575 2.805 ;
        RECT 14.865 2.635 15.035 2.805 ;
        RECT 15.325 2.635 15.495 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
        RECT 14.405 -0.085 14.575 0.085 ;
        RECT 14.865 -0.085 15.035 0.085 ;
        RECT 15.325 -0.085 15.495 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand2_16

#--------EOF---------

MACRO sky130_fd_sc_hdll__nand2b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand2b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 0.420 1.315 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.590 1.075 1.185 1.315 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.335 1.990 1.015 ;
        RECT 0.150 0.105 1.990 0.335 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.491500 ;
    PORT
      LAYER li1 ;
        RECT 1.050 2.005 1.430 2.465 ;
        RECT 1.050 1.835 2.190 2.005 ;
        RECT 1.820 0.545 2.190 1.835 ;
        RECT 1.360 0.255 2.190 0.545 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.630 1.835 0.880 2.635 ;
        RECT 1.650 2.175 1.865 2.635 ;
        RECT 0.090 1.665 0.370 1.825 ;
        RECT 0.090 1.495 1.620 1.665 ;
        RECT 1.450 0.905 1.620 1.495 ;
        RECT 0.090 0.735 1.620 0.905 ;
        RECT 0.090 0.525 0.360 0.735 ;
        RECT 0.630 0.085 0.960 0.545 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand2b_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__nand2b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand2b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.455 0.995 0.850 1.325 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.905 1.275 3.095 1.655 ;
        RECT 2.110 1.075 3.095 1.275 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.335 3.185 1.015 ;
        RECT 0.150 0.105 3.185 0.335 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.825500 ;
    PORT
      LAYER li1 ;
        RECT 1.135 2.005 1.465 2.465 ;
        RECT 2.285 2.005 2.615 2.465 ;
        RECT 1.135 1.835 2.615 2.005 ;
        RECT 1.455 0.635 1.785 1.835 ;
        RECT 2.340 1.495 2.615 1.835 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.110 1.665 0.410 1.860 ;
        RECT 0.630 1.835 0.885 2.635 ;
        RECT 1.725 2.175 2.100 2.635 ;
        RECT 2.845 1.835 3.015 2.635 ;
        RECT 0.110 1.495 1.190 1.665 ;
        RECT 0.110 0.840 0.280 1.495 ;
        RECT 1.020 0.995 1.190 1.495 ;
        RECT 0.110 0.510 0.345 0.840 ;
        RECT 0.595 0.085 0.765 0.775 ;
        RECT 1.955 0.695 3.095 0.905 ;
        RECT 1.955 0.465 2.205 0.695 ;
        RECT 1.035 0.255 2.205 0.465 ;
        RECT 2.425 0.085 2.595 0.525 ;
        RECT 2.765 0.255 3.095 0.695 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand2b_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__nand2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand2b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.110 1.075 0.440 1.275 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 3.405 1.075 5.390 1.275 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.410 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.576000 ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.665 1.885 2.465 ;
        RECT 2.445 1.665 2.840 2.465 ;
        RECT 3.400 1.665 3.780 2.465 ;
        RECT 4.340 1.665 4.720 2.465 ;
        RECT 1.505 1.445 4.720 1.665 ;
        RECT 2.575 0.905 2.840 1.445 ;
        RECT 1.505 0.635 2.840 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.090 1.665 0.425 2.465 ;
        RECT 0.645 1.835 1.335 2.635 ;
        RECT 2.105 1.835 2.275 2.635 ;
        RECT 3.060 1.835 3.230 2.635 ;
        RECT 4.000 1.835 4.170 2.635 ;
        RECT 0.090 1.445 0.830 1.665 ;
        RECT 1.020 1.445 1.335 1.835 ;
        RECT 4.970 1.495 5.300 2.635 ;
        RECT 0.660 1.275 0.830 1.445 ;
        RECT 0.660 1.075 2.355 1.275 ;
        RECT 0.660 0.905 0.830 1.075 ;
        RECT 0.090 0.715 0.830 0.905 ;
        RECT 0.090 0.255 0.425 0.715 ;
        RECT 0.645 0.085 0.840 0.545 ;
        RECT 1.085 0.465 1.335 0.905 ;
        RECT 3.060 0.715 5.300 0.905 ;
        RECT 3.060 0.465 3.310 0.715 ;
        RECT 1.085 0.255 3.310 0.465 ;
        RECT 3.530 0.085 3.700 0.545 ;
        RECT 3.870 0.255 4.250 0.715 ;
        RECT 4.470 0.085 4.710 0.545 ;
        RECT 4.970 0.255 5.300 0.715 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand2b_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__nand3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.475 0.995 1.905 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.915 0.765 1.285 1.325 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.110 0.745 0.330 1.325 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 1.985 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.761500 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.665 0.895 2.465 ;
        RECT 1.515 1.665 1.895 2.465 ;
        RECT 0.515 1.495 1.895 1.665 ;
        RECT 0.515 0.595 0.745 1.495 ;
        RECT 1.515 0.595 1.895 0.825 ;
        RECT 0.515 0.255 1.895 0.595 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.090 1.495 0.345 2.635 ;
        RECT 1.115 1.835 1.345 2.635 ;
        RECT 0.090 0.085 0.345 0.575 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand3_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__nand3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.995 0.330 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 1.170 1.075 2.615 1.275 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.785 1.075 4.000 1.275 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.905 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.078000 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.665 0.895 2.465 ;
        RECT 1.455 1.665 1.835 2.465 ;
        RECT 2.915 1.665 3.295 2.465 ;
        RECT 0.515 1.445 3.295 1.665 ;
        RECT 0.515 0.635 0.895 1.445 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.090 1.495 0.345 2.635 ;
        RECT 1.115 1.835 1.285 2.635 ;
        RECT 2.055 1.835 2.745 2.635 ;
        RECT 3.515 1.445 3.895 2.635 ;
        RECT 0.090 0.465 0.345 0.785 ;
        RECT 1.455 0.635 3.295 0.905 ;
        RECT 0.090 0.295 2.305 0.465 ;
        RECT 2.495 0.085 2.825 0.465 ;
        RECT 3.515 0.085 3.895 0.885 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand3_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__nand3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.900 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 4.250 1.075 6.370 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 2.275 1.075 4.025 1.275 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.110 1.075 1.850 1.275 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.900 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 6.685 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.090 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.900 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.156000 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.665 0.895 2.465 ;
        RECT 1.455 1.665 1.835 2.465 ;
        RECT 2.395 1.665 2.775 2.465 ;
        RECT 3.335 1.665 3.715 2.465 ;
        RECT 4.795 1.665 5.175 2.465 ;
        RECT 5.735 1.665 6.115 2.465 ;
        RECT 0.515 1.445 6.785 1.665 ;
        RECT 6.555 0.905 6.785 1.445 ;
        RECT 4.795 0.655 6.785 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.900 2.805 ;
        RECT 0.090 1.445 0.345 2.635 ;
        RECT 1.115 1.835 1.285 2.635 ;
        RECT 2.055 1.835 2.225 2.635 ;
        RECT 2.995 1.835 3.165 2.635 ;
        RECT 3.935 1.835 4.625 2.635 ;
        RECT 5.395 1.835 5.565 2.635 ;
        RECT 6.335 1.835 6.600 2.635 ;
        RECT 0.090 0.735 4.185 0.905 ;
        RECT 0.090 0.255 0.425 0.735 ;
        RECT 0.645 0.085 0.815 0.565 ;
        RECT 0.985 0.255 1.365 0.735 ;
        RECT 1.925 0.655 2.305 0.735 ;
        RECT 2.865 0.655 3.245 0.735 ;
        RECT 3.805 0.655 4.185 0.735 ;
        RECT 1.585 0.085 1.755 0.565 ;
        RECT 2.395 0.255 6.600 0.485 ;
        RECT 0.000 -0.085 6.900 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand3_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__nand3b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand3b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.995 0.825 1.325 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.520 0.995 1.795 1.325 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.015 0.995 1.335 1.325 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.135 0.335 2.630 1.015 ;
        RECT 0.145 0.105 2.630 0.335 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.775250 ;
    PORT
      LAYER li1 ;
        RECT 1.180 1.665 1.560 2.465 ;
        RECT 2.130 1.665 2.675 2.465 ;
        RECT 1.180 1.495 2.675 1.665 ;
        RECT 2.410 0.485 2.675 1.495 ;
        RECT 2.130 0.255 2.675 0.485 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.085 1.595 0.510 1.925 ;
        RECT 0.085 0.825 0.255 1.595 ;
        RECT 0.760 1.495 1.010 2.635 ;
        RECT 1.790 1.835 1.960 2.635 ;
        RECT 2.000 0.825 2.220 1.325 ;
        RECT 0.085 0.655 2.220 0.825 ;
        RECT 0.085 0.445 0.510 0.655 ;
        RECT 0.760 0.085 1.090 0.485 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand3b_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__nand3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand3b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.430 1.075 0.830 1.275 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.150 1.075 3.440 1.275 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.075 1.890 1.275 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.540 0.785 4.500 1.015 ;
        RECT 0.005 0.105 4.500 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.110500 ;
    PORT
      LAYER li1 ;
        RECT 1.110 2.005 1.490 2.465 ;
        RECT 2.050 2.005 2.430 2.465 ;
        RECT 1.110 1.955 2.430 2.005 ;
        RECT 3.560 2.005 3.860 2.465 ;
        RECT 3.560 1.955 4.490 2.005 ;
        RECT 1.110 1.785 4.490 1.955 ;
        RECT 4.250 0.905 4.490 1.785 ;
        RECT 3.560 0.635 4.490 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.090 2.065 0.410 2.465 ;
        RECT 0.090 1.615 0.260 2.065 ;
        RECT 0.630 1.835 0.940 2.635 ;
        RECT 1.710 2.175 1.880 2.635 ;
        RECT 2.650 2.175 2.900 2.635 ;
        RECT 3.090 2.175 3.390 2.635 ;
        RECT 4.160 2.175 4.450 2.635 ;
        RECT 0.090 1.445 4.000 1.615 ;
        RECT 0.090 0.655 0.260 1.445 ;
        RECT 3.670 1.075 4.000 1.445 ;
        RECT 0.090 0.255 0.410 0.655 ;
        RECT 0.630 0.085 0.940 0.905 ;
        RECT 1.110 0.715 3.000 0.905 ;
        RECT 1.110 0.255 1.490 0.715 ;
        RECT 2.200 0.635 3.000 0.715 ;
        RECT 1.710 0.085 1.960 0.545 ;
        RECT 3.220 0.465 3.390 0.905 ;
        RECT 2.200 0.255 4.450 0.465 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand3b_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__nand3b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand3b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.820 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.430 1.075 0.830 1.275 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 3.725 1.075 4.930 1.275 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 5.185 1.075 7.100 1.275 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.820 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 7.765 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.010 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.820 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.156000 ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.665 1.885 2.465 ;
        RECT 2.445 2.005 2.825 2.465 ;
        RECT 3.385 2.005 3.765 2.465 ;
        RECT 2.445 1.665 3.765 2.005 ;
        RECT 4.325 1.665 4.705 2.465 ;
        RECT 5.785 1.665 6.165 2.465 ;
        RECT 6.725 1.665 7.105 2.465 ;
        RECT 1.505 1.445 7.105 1.665 ;
        RECT 3.045 1.075 3.555 1.445 ;
        RECT 3.045 0.905 3.215 1.075 ;
        RECT 1.505 0.635 3.215 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.820 2.805 ;
        RECT 0.085 1.445 0.425 2.465 ;
        RECT 0.645 1.445 1.335 2.635 ;
        RECT 2.105 1.835 2.275 2.635 ;
        RECT 3.045 2.175 3.215 2.635 ;
        RECT 3.985 1.835 4.155 2.635 ;
        RECT 4.925 1.835 5.615 2.635 ;
        RECT 6.385 1.835 6.555 2.635 ;
        RECT 7.325 1.445 7.655 2.635 ;
        RECT 0.085 0.905 0.260 1.445 ;
        RECT 1.055 1.075 2.825 1.275 ;
        RECT 1.055 0.905 1.335 1.075 ;
        RECT 0.085 0.715 1.335 0.905 ;
        RECT 3.385 0.715 7.105 0.905 ;
        RECT 0.085 0.255 0.425 0.715 ;
        RECT 3.385 0.635 5.175 0.715 ;
        RECT 0.645 0.085 0.895 0.545 ;
        RECT 1.085 0.255 5.175 0.465 ;
        RECT 5.365 0.085 5.615 0.545 ;
        RECT 5.785 0.255 6.165 0.715 ;
        RECT 6.385 0.085 6.555 0.545 ;
        RECT 6.725 0.255 7.105 0.715 ;
        RECT 7.325 0.085 7.655 0.905 ;
        RECT 0.000 -0.085 7.820 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand3b_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__nand4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.175 0.995 2.640 1.665 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.245 0.995 1.605 1.325 ;
        RECT 1.245 0.825 1.415 0.995 ;
        RECT 1.030 0.300 1.415 0.825 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.595 0.995 1.075 1.325 ;
        RECT 0.595 0.300 0.860 0.995 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.110 0.995 0.395 1.325 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.495 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.867500 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.665 0.895 2.465 ;
        RECT 1.535 1.665 1.865 2.465 ;
        RECT 0.515 1.495 1.945 1.665 ;
        RECT 1.775 0.825 1.945 1.495 ;
        RECT 1.670 0.255 2.415 0.825 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.085 1.495 0.345 2.635 ;
        RECT 1.115 1.835 1.285 2.635 ;
        RECT 2.115 1.835 2.395 2.635 ;
        RECT 0.090 0.085 0.425 0.825 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand4_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__nand4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 4.615 1.075 4.945 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.435 1.075 3.380 1.275 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.075 1.850 1.275 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.110 1.075 0.895 1.275 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.985 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.368000 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.665 0.895 2.465 ;
        RECT 1.455 1.665 1.835 2.465 ;
        RECT 2.555 1.665 2.935 2.465 ;
        RECT 3.945 1.665 4.325 2.465 ;
        RECT 0.515 1.445 4.325 1.665 ;
        RECT 3.720 1.055 4.325 1.445 ;
        RECT 3.945 0.635 4.325 1.055 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.060 2.805 ;
        RECT 0.090 1.495 0.345 2.635 ;
        RECT 1.115 1.835 1.285 2.635 ;
        RECT 2.055 1.835 2.385 2.635 ;
        RECT 3.295 1.835 3.675 2.635 ;
        RECT 4.545 1.445 4.875 2.635 ;
        RECT 0.090 0.735 1.285 0.905 ;
        RECT 0.090 0.255 0.425 0.735 ;
        RECT 0.645 0.085 0.815 0.545 ;
        RECT 0.985 0.465 1.285 0.735 ;
        RECT 1.455 0.635 3.385 0.905 ;
        RECT 3.605 0.465 3.775 0.885 ;
        RECT 4.545 0.465 4.875 0.905 ;
        RECT 0.985 0.255 2.325 0.465 ;
        RECT 2.515 0.255 4.875 0.465 ;
        RECT 0.000 -0.085 5.060 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand4_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__nand4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.740 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 7.115 1.075 8.510 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 4.250 1.075 6.115 1.275 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 2.190 1.075 4.025 1.275 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 1.835 1.275 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.740 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 8.615 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.925 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.740 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.736000 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.665 0.895 2.465 ;
        RECT 1.455 1.665 1.835 2.465 ;
        RECT 2.395 1.665 2.775 2.465 ;
        RECT 3.335 1.665 3.715 2.465 ;
        RECT 4.795 1.665 5.175 2.465 ;
        RECT 5.735 1.665 6.115 2.465 ;
        RECT 6.735 1.665 7.115 2.465 ;
        RECT 7.675 1.665 8.055 2.465 ;
        RECT 0.515 1.445 8.055 1.665 ;
        RECT 6.545 0.905 6.825 1.445 ;
        RECT 6.545 0.655 8.055 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.740 2.805 ;
        RECT 0.090 1.445 0.345 2.635 ;
        RECT 1.115 1.835 1.285 2.635 ;
        RECT 2.055 1.835 2.225 2.635 ;
        RECT 2.995 1.835 3.165 2.635 ;
        RECT 3.935 1.835 4.625 2.635 ;
        RECT 5.395 1.835 5.565 2.635 ;
        RECT 6.370 1.835 6.540 2.635 ;
        RECT 7.335 1.835 7.505 2.635 ;
        RECT 8.275 1.445 8.535 2.635 ;
        RECT 0.090 0.655 2.225 0.905 ;
        RECT 2.395 0.655 6.115 0.905 ;
        RECT 0.090 0.255 0.345 0.655 ;
        RECT 0.515 0.085 0.895 0.485 ;
        RECT 1.115 0.255 1.285 0.655 ;
        RECT 2.055 0.485 2.225 0.655 ;
        RECT 8.275 0.485 8.530 0.905 ;
        RECT 1.455 0.085 1.835 0.485 ;
        RECT 2.055 0.255 4.185 0.485 ;
        RECT 4.375 0.255 8.530 0.485 ;
        RECT 0.000 -0.085 8.740 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand4_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__nand4b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand4b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.995 0.820 1.325 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.930 0.765 2.225 1.325 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.500 0.960 1.760 1.325 ;
        RECT 1.540 0.765 1.760 0.960 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.010 0.995 1.330 1.325 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.070 0.335 3.215 1.015 ;
        RECT 0.145 0.105 3.215 0.335 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.882500 ;
    PORT
      LAYER li1 ;
        RECT 1.175 1.665 1.555 2.465 ;
        RECT 2.175 1.665 2.505 2.465 ;
        RECT 1.175 1.495 3.135 1.665 ;
        RECT 2.875 0.835 3.135 1.495 ;
        RECT 2.775 0.255 3.135 0.835 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.085 1.595 0.505 1.925 ;
        RECT 0.085 0.825 0.255 1.595 ;
        RECT 0.755 1.495 1.005 2.635 ;
        RECT 1.725 1.835 2.000 2.635 ;
        RECT 2.875 1.835 3.090 2.635 ;
        RECT 2.395 0.995 2.705 1.325 ;
        RECT 0.085 0.655 1.370 0.825 ;
        RECT 0.085 0.445 0.470 0.655 ;
        RECT 1.200 0.595 1.370 0.655 ;
        RECT 2.395 0.595 2.600 0.995 ;
        RECT 0.665 0.085 1.030 0.485 ;
        RECT 1.200 0.425 2.600 0.595 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand4b_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__nand4b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand4b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.995 0.330 1.615 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.160 1.075 3.350 1.275 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 3.610 1.075 4.685 1.275 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 5.020 1.075 5.885 1.275 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.995 0.785 5.875 1.015 ;
        RECT 0.005 0.105 5.875 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.368000 ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.665 1.885 2.465 ;
        RECT 2.445 1.665 2.825 2.465 ;
        RECT 3.855 1.665 4.235 2.465 ;
        RECT 4.885 1.665 5.265 2.465 ;
        RECT 1.505 1.445 5.265 1.665 ;
        RECT 1.505 0.635 1.885 1.445 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.090 2.085 0.345 2.465 ;
        RECT 0.515 2.255 1.335 2.635 ;
        RECT 0.090 1.915 0.720 2.085 ;
        RECT 0.500 1.245 0.720 1.915 ;
        RECT 1.085 1.445 1.335 2.255 ;
        RECT 2.105 1.835 2.275 2.635 ;
        RECT 3.045 1.835 3.685 2.635 ;
        RECT 4.455 1.835 4.715 2.635 ;
        RECT 5.485 1.495 5.880 2.635 ;
        RECT 0.500 1.075 1.335 1.245 ;
        RECT 0.500 0.805 0.720 1.075 ;
        RECT 0.090 0.635 0.720 0.805 ;
        RECT 0.090 0.255 0.345 0.635 ;
        RECT 1.085 0.465 1.335 0.905 ;
        RECT 2.105 0.635 3.295 0.905 ;
        RECT 3.485 0.715 5.790 0.905 ;
        RECT 3.485 0.635 4.805 0.715 ;
        RECT 2.105 0.465 2.275 0.635 ;
        RECT 4.505 0.615 4.805 0.635 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.085 0.255 2.275 0.465 ;
        RECT 2.445 0.255 4.285 0.465 ;
        RECT 4.505 0.255 4.765 0.615 ;
        RECT 5.065 0.085 5.235 0.545 ;
        RECT 5.455 0.255 5.790 0.715 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand4b_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__nand4b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand4b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.660 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.110 1.075 0.440 1.275 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 3.180 1.075 5.040 1.275 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 5.240 1.075 7.110 1.275 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 7.665 1.075 9.505 1.275 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.660 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 9.545 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.850 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.660 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.736000 ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.665 1.885 2.465 ;
        RECT 2.445 1.665 2.825 2.465 ;
        RECT 3.385 1.665 3.765 2.465 ;
        RECT 4.325 1.665 4.705 2.465 ;
        RECT 5.785 1.665 6.165 2.465 ;
        RECT 6.725 1.665 7.105 2.465 ;
        RECT 7.665 1.665 8.045 2.465 ;
        RECT 8.605 1.665 8.985 2.465 ;
        RECT 1.505 1.445 8.985 1.665 ;
        RECT 2.410 0.905 2.840 1.445 ;
        RECT 1.505 0.635 2.840 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.660 2.805 ;
        RECT 0.090 1.665 0.425 2.465 ;
        RECT 0.645 1.835 1.335 2.635 ;
        RECT 2.105 1.835 2.275 2.635 ;
        RECT 3.045 1.835 3.215 2.635 ;
        RECT 3.985 1.835 4.155 2.635 ;
        RECT 4.925 1.835 5.615 2.635 ;
        RECT 6.385 1.835 6.555 2.635 ;
        RECT 7.325 1.835 7.495 2.635 ;
        RECT 8.265 1.835 8.435 2.635 ;
        RECT 0.090 1.495 0.855 1.665 ;
        RECT 1.045 1.495 1.335 1.835 ;
        RECT 0.660 1.275 0.855 1.495 ;
        RECT 9.205 1.445 9.460 2.635 ;
        RECT 0.660 1.075 1.975 1.275 ;
        RECT 0.660 0.905 0.855 1.075 ;
        RECT 0.090 0.735 0.855 0.905 ;
        RECT 0.090 0.255 0.425 0.735 ;
        RECT 0.645 0.085 0.895 0.545 ;
        RECT 1.085 0.465 1.335 0.905 ;
        RECT 3.385 0.635 7.105 0.905 ;
        RECT 7.325 0.735 9.460 0.905 ;
        RECT 7.325 0.465 7.575 0.735 ;
        RECT 1.085 0.255 5.175 0.465 ;
        RECT 5.365 0.255 7.575 0.465 ;
        RECT 7.795 0.085 7.965 0.545 ;
        RECT 8.135 0.255 8.515 0.735 ;
        RECT 8.735 0.085 8.905 0.545 ;
        RECT 9.075 0.255 9.460 0.735 ;
        RECT 0.000 -0.085 9.660 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand4b_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__nand4bb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand4bb_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 3.300 0.725 3.710 1.615 ;
    END
  END A_N
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.430 1.075 0.825 1.655 ;
    END
  END B_N
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.495 0.735 1.760 1.325 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.995 1.075 1.325 1.325 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.785 3.090 1.015 ;
        RECT 0.005 0.335 4.135 0.785 ;
        RECT 0.145 0.105 4.135 0.335 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.901500 ;
    PORT
      LAYER li1 ;
        RECT 1.155 1.665 1.485 2.465 ;
        RECT 2.190 2.005 2.580 2.465 ;
        RECT 2.190 1.665 2.680 2.005 ;
        RECT 1.155 1.495 2.680 1.665 ;
        RECT 2.410 0.825 2.680 1.495 ;
        RECT 2.410 0.255 3.000 0.825 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.085 2.065 0.425 2.465 ;
        RECT 0.085 0.905 0.260 2.065 ;
        RECT 0.645 1.835 0.975 2.635 ;
        RECT 1.695 1.835 2.015 2.635 ;
        RECT 2.750 2.175 3.520 2.635 ;
        RECT 3.740 2.005 4.055 2.465 ;
        RECT 2.850 1.835 4.055 2.005 ;
        RECT 0.085 0.715 1.220 0.905 ;
        RECT 0.085 0.485 0.425 0.715 ;
        RECT 1.050 0.555 1.220 0.715 ;
        RECT 1.990 0.555 2.240 1.325 ;
        RECT 2.850 0.995 3.125 1.835 ;
        RECT 0.645 0.085 0.880 0.545 ;
        RECT 1.050 0.365 2.240 0.555 ;
        RECT 3.885 0.545 4.055 1.835 ;
        RECT 3.190 0.085 3.540 0.545 ;
        RECT 3.710 0.255 4.055 0.545 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand4bb_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__nand4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand4bb_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.560 1.070 0.940 1.615 ;
    END
  END A_N
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.070 0.330 1.615 ;
    END
  END B_N
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 4.240 1.075 4.950 1.275 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 5.315 1.075 6.295 1.275 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.675 0.785 6.435 1.015 ;
        RECT 0.005 0.105 6.435 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.368000 ;
    PORT
      LAYER li1 ;
        RECT 2.185 1.665 2.485 2.465 ;
        RECT 3.125 1.665 3.505 2.465 ;
        RECT 4.555 1.665 4.935 2.465 ;
        RECT 5.495 1.665 5.875 2.465 ;
        RECT 2.185 1.445 5.875 1.665 ;
        RECT 2.185 0.655 2.630 1.445 ;
        RECT 3.495 1.075 4.045 1.445 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.085 1.980 0.370 2.440 ;
        RECT 0.540 2.195 0.815 2.635 ;
        RECT 0.985 2.150 1.675 2.465 ;
        RECT 0.085 1.785 1.330 1.980 ;
        RECT 1.160 0.900 1.330 1.785 ;
        RECT 0.085 0.730 1.330 0.900 ;
        RECT 0.085 0.255 0.345 0.730 ;
        RECT 1.500 0.560 1.675 2.150 ;
        RECT 1.845 1.495 2.015 2.635 ;
        RECT 2.655 1.835 2.955 2.635 ;
        RECT 3.725 1.835 4.385 2.635 ;
        RECT 5.155 1.835 5.325 2.635 ;
        RECT 6.095 1.445 6.345 2.635 ;
        RECT 2.945 1.075 3.325 1.275 ;
        RECT 3.125 0.655 4.935 0.905 ;
        RECT 5.155 0.735 6.345 0.905 ;
        RECT 0.515 0.085 0.815 0.545 ;
        RECT 0.985 0.255 1.675 0.560 ;
        RECT 1.845 0.485 2.015 0.585 ;
        RECT 5.155 0.485 5.405 0.735 ;
        RECT 1.845 0.255 3.975 0.485 ;
        RECT 4.165 0.255 5.405 0.485 ;
        RECT 5.625 0.085 5.795 0.565 ;
        RECT 5.965 0.255 6.345 0.735 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 1.160 1.105 1.330 1.275 ;
        RECT 3.155 1.105 3.325 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
      LAYER met1 ;
        RECT 1.100 1.075 3.385 1.305 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand4bb_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__nand4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand4bb_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.580 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.100 0.995 0.330 1.615 ;
    END
  END A_N
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.585 0.995 1.025 1.615 ;
    END
  END B_N
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 6.045 1.075 7.985 1.275 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 8.395 1.075 10.340 1.275 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.580 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 10.440 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.770 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.580 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.736000 ;
    PORT
      LAYER li1 ;
        RECT 2.355 1.665 2.655 2.465 ;
        RECT 3.295 1.665 3.675 2.465 ;
        RECT 4.235 1.665 4.615 2.465 ;
        RECT 5.175 1.665 5.555 2.465 ;
        RECT 6.665 1.665 7.045 2.465 ;
        RECT 7.605 1.665 7.985 2.465 ;
        RECT 8.545 1.665 8.925 2.465 ;
        RECT 9.485 1.665 9.865 2.465 ;
        RECT 2.355 1.445 9.865 1.665 ;
        RECT 3.665 0.905 4.015 1.445 ;
        RECT 2.355 0.655 4.015 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.580 2.805 ;
        RECT 0.085 1.980 0.370 2.440 ;
        RECT 0.540 2.195 0.815 2.635 ;
        RECT 0.985 2.150 1.845 2.465 ;
        RECT 0.085 1.785 1.505 1.980 ;
        RECT 1.195 0.805 1.505 1.785 ;
        RECT 0.085 0.635 1.505 0.805 ;
        RECT 1.675 1.305 1.845 2.150 ;
        RECT 2.015 1.495 2.185 2.635 ;
        RECT 2.825 1.835 3.125 2.635 ;
        RECT 3.895 1.835 4.065 2.635 ;
        RECT 4.835 1.835 5.005 2.635 ;
        RECT 5.825 1.835 6.465 2.635 ;
        RECT 7.265 1.835 7.435 2.635 ;
        RECT 8.205 1.835 8.375 2.635 ;
        RECT 9.145 1.835 9.315 2.635 ;
        RECT 10.085 1.445 10.360 2.635 ;
        RECT 1.675 1.075 2.025 1.305 ;
        RECT 2.355 1.075 3.200 1.245 ;
        RECT 4.185 1.075 5.555 1.275 ;
        RECT 0.085 0.255 0.345 0.635 ;
        RECT 1.675 0.465 1.845 1.075 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.115 0.255 1.845 0.465 ;
        RECT 2.015 0.485 2.185 0.905 ;
        RECT 4.235 0.655 8.010 0.905 ;
        RECT 8.205 0.655 10.285 0.825 ;
        RECT 8.205 0.485 8.375 0.655 ;
        RECT 2.015 0.255 6.025 0.485 ;
        RECT 6.265 0.255 8.375 0.485 ;
        RECT 8.595 0.085 8.925 0.485 ;
        RECT 9.535 0.085 9.865 0.485 ;
        RECT 0.000 -0.085 10.580 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 1.795 1.105 1.965 1.275 ;
        RECT 4.330 1.105 4.500 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
      LAYER met1 ;
        RECT 1.735 1.260 2.025 1.305 ;
        RECT 4.235 1.260 4.575 1.305 ;
        RECT 1.735 1.120 4.575 1.260 ;
        RECT 1.735 1.075 2.025 1.120 ;
        RECT 4.235 1.075 4.575 1.120 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand4bb_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__nor2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nor2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.045 1.075 1.395 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.435 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 1.745 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.665 0.425 2.450 ;
        RECT 0.095 1.495 0.775 1.665 ;
        RECT 0.605 0.895 0.775 1.495 ;
        RECT 0.515 0.255 0.895 0.895 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.840 2.805 ;
        RECT 1.115 1.495 1.625 2.635 ;
        RECT 0.105 0.085 0.345 0.895 ;
        RECT 1.065 0.085 1.575 0.895 ;
        RECT 0.000 -0.085 1.840 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor2_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__nor2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nor2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 0.860 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 1.030 1.075 1.900 1.275 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.530 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.771000 ;
    PORT
      LAYER li1 ;
        RECT 1.475 1.665 1.855 2.125 ;
        RECT 1.475 1.445 2.310 1.665 ;
        RECT 2.095 0.905 2.310 1.445 ;
        RECT 0.535 0.735 2.310 0.905 ;
        RECT 0.535 0.725 1.855 0.735 ;
        RECT 0.535 0.255 0.915 0.725 ;
        RECT 1.475 0.255 1.855 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.090 1.665 0.365 2.465 ;
        RECT 0.535 1.835 0.915 2.635 ;
        RECT 1.135 2.295 2.375 2.465 ;
        RECT 1.135 1.665 1.305 2.295 ;
        RECT 2.075 1.835 2.375 2.295 ;
        RECT 0.090 1.455 1.305 1.665 ;
        RECT 0.090 0.085 0.365 0.905 ;
        RECT 1.135 0.085 1.305 0.555 ;
        RECT 2.140 0.085 2.480 0.555 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor2_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__nor2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nor2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.140 1.075 1.950 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 2.320 1.075 3.835 1.275 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.295 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.477000 ;
    PORT
      LAYER li1 ;
        RECT 2.545 1.745 2.715 2.125 ;
        RECT 3.485 1.745 3.655 2.125 ;
        RECT 2.545 1.445 4.490 1.745 ;
        RECT 4.095 0.905 4.490 1.445 ;
        RECT 0.535 0.725 4.490 0.905 ;
        RECT 0.535 0.255 0.915 0.725 ;
        RECT 1.475 0.255 1.855 0.725 ;
        RECT 2.415 0.255 2.795 0.725 ;
        RECT 3.355 0.255 3.735 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.090 1.665 0.365 2.465 ;
        RECT 0.535 1.835 0.915 2.635 ;
        RECT 1.135 1.665 1.305 2.465 ;
        RECT 1.475 1.835 1.775 2.635 ;
        RECT 1.945 2.295 4.290 2.465 ;
        RECT 1.945 1.665 2.325 2.295 ;
        RECT 2.885 1.935 3.265 2.295 ;
        RECT 3.825 1.915 4.290 2.295 ;
        RECT 0.090 1.455 2.325 1.665 ;
        RECT 0.090 0.085 0.365 0.905 ;
        RECT 1.135 0.085 1.305 0.555 ;
        RECT 2.075 0.085 2.245 0.555 ;
        RECT 3.015 0.085 3.185 0.555 ;
        RECT 3.955 0.085 4.240 0.555 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor2_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__nor2_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nor2_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.280 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.220000 ;
    PORT
      LAYER li1 ;
        RECT 0.360 1.075 3.930 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.220000 ;
    PORT
      LAYER li1 ;
        RECT 4.200 1.075 7.290 1.275 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.280 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 8.055 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.470 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.280 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.889000 ;
    PORT
      LAYER li1 ;
        RECT 4.385 1.615 4.635 2.125 ;
        RECT 5.325 1.615 5.575 2.125 ;
        RECT 6.265 1.615 6.515 2.125 ;
        RECT 7.205 1.615 7.455 2.125 ;
        RECT 4.385 1.445 8.025 1.615 ;
        RECT 7.460 0.905 8.025 1.445 ;
        RECT 0.535 0.725 8.025 0.905 ;
        RECT 0.535 0.255 0.915 0.725 ;
        RECT 1.475 0.255 1.855 0.725 ;
        RECT 2.415 0.255 2.795 0.725 ;
        RECT 3.355 0.255 3.735 0.725 ;
        RECT 4.295 0.255 4.675 0.725 ;
        RECT 5.235 0.255 5.615 0.725 ;
        RECT 6.175 0.255 6.555 0.725 ;
        RECT 7.115 0.255 7.495 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.280 2.805 ;
        RECT 0.090 1.665 0.405 2.465 ;
        RECT 0.625 1.835 0.875 2.635 ;
        RECT 1.095 1.665 1.345 2.465 ;
        RECT 1.565 1.835 1.815 2.635 ;
        RECT 2.035 1.665 2.285 2.465 ;
        RECT 2.505 1.835 2.755 2.635 ;
        RECT 2.975 1.665 3.225 2.465 ;
        RECT 3.445 1.835 3.695 2.635 ;
        RECT 3.915 2.295 7.925 2.465 ;
        RECT 3.915 1.665 4.165 2.295 ;
        RECT 4.855 1.785 5.105 2.295 ;
        RECT 5.795 1.785 6.045 2.295 ;
        RECT 6.735 1.785 6.985 2.295 ;
        RECT 7.675 1.785 7.925 2.295 ;
        RECT 0.090 1.455 4.165 1.665 ;
        RECT 0.090 0.085 0.365 0.905 ;
        RECT 1.135 0.085 1.305 0.555 ;
        RECT 2.075 0.085 2.245 0.555 ;
        RECT 3.015 0.085 3.185 0.555 ;
        RECT 3.955 0.085 4.125 0.555 ;
        RECT 4.895 0.085 5.065 0.555 ;
        RECT 5.835 0.085 6.005 0.555 ;
        RECT 6.775 0.085 6.945 0.555 ;
        RECT 7.715 0.085 8.005 0.555 ;
        RECT 0.000 -0.085 8.280 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor2_8

#--------EOF---------

MACRO sky130_fd_sc_hdll__nor2b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nor2b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.955 1.065 1.285 1.325 ;
    END
  END A
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.975 0.785 1.745 ;
    END
  END B_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.625 0.785 2.075 1.015 ;
        RECT 0.005 0.105 2.075 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 1.655 1.850 2.215 2.465 ;
        RECT 2.035 0.895 2.215 1.850 ;
        RECT 1.135 0.725 2.215 0.895 ;
        RECT 1.135 0.255 1.515 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.775 2.255 1.105 2.635 ;
        RECT 0.095 1.915 1.485 2.085 ;
        RECT 0.095 0.290 0.345 1.915 ;
        RECT 1.315 1.665 1.485 1.915 ;
        RECT 1.315 1.495 1.655 1.665 ;
        RECT 1.485 1.325 1.655 1.495 ;
        RECT 1.485 1.075 1.865 1.325 ;
        RECT 0.675 0.085 0.965 0.625 ;
        RECT 1.735 0.085 2.120 0.555 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor2b_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__nor2b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nor2b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.480 1.065 1.260 1.275 ;
    END
  END A
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 3.270 1.275 3.535 1.965 ;
        RECT 2.960 1.065 3.535 1.275 ;
    END
  END B_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.335 3.565 1.015 ;
        RECT 0.010 0.105 2.415 0.335 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.738500 ;
    PORT
      LAYER li1 ;
        RECT 1.565 0.895 1.815 2.125 ;
        RECT 0.535 0.725 1.855 0.895 ;
        RECT 0.535 0.255 0.935 0.725 ;
        RECT 1.475 0.255 1.855 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.085 1.655 0.405 2.465 ;
        RECT 0.625 1.825 0.875 2.635 ;
        RECT 1.095 2.295 2.325 2.465 ;
        RECT 1.095 1.655 1.345 2.295 ;
        RECT 0.085 1.445 1.345 1.655 ;
        RECT 2.035 1.445 2.325 2.295 ;
        RECT 2.595 1.245 2.765 2.460 ;
        RECT 3.185 2.145 3.435 2.635 ;
        RECT 2.075 1.075 2.765 1.245 ;
        RECT 0.085 0.085 0.365 0.895 ;
        RECT 1.135 0.085 1.305 0.555 ;
        RECT 2.075 0.085 2.245 0.895 ;
        RECT 2.595 0.445 2.765 1.075 ;
        RECT 3.185 0.085 3.440 0.845 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor2b_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__nor2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nor2b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.360 1.075 1.950 1.275 ;
    END
  END A
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.075 5.425 1.320 ;
    END
  END B_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.325 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444500 ;
    PORT
      LAYER li1 ;
        RECT 2.545 1.745 2.715 2.125 ;
        RECT 3.485 1.745 3.655 2.125 ;
        RECT 2.545 1.415 3.655 1.745 ;
        RECT 2.545 0.905 2.875 1.415 ;
        RECT 0.535 0.725 3.735 0.905 ;
        RECT 0.535 0.255 0.915 0.725 ;
        RECT 1.475 0.255 1.855 0.725 ;
        RECT 2.415 0.255 2.795 0.725 ;
        RECT 3.355 0.255 3.735 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.085 1.665 0.365 2.465 ;
        RECT 0.535 1.835 0.915 2.635 ;
        RECT 1.135 1.665 1.305 2.465 ;
        RECT 1.475 1.835 1.775 2.635 ;
        RECT 1.945 2.295 4.225 2.465 ;
        RECT 1.945 1.665 2.325 2.295 ;
        RECT 2.885 1.935 3.265 2.295 ;
        RECT 0.085 1.455 2.325 1.665 ;
        RECT 3.825 1.575 4.225 2.295 ;
        RECT 4.395 1.245 4.755 2.465 ;
        RECT 4.975 1.495 5.380 2.635 ;
        RECT 3.065 1.075 4.755 1.245 ;
        RECT 0.085 0.085 0.365 0.905 ;
        RECT 1.135 0.085 1.305 0.555 ;
        RECT 2.075 0.085 2.245 0.555 ;
        RECT 3.015 0.085 3.185 0.555 ;
        RECT 3.955 0.085 4.125 0.905 ;
        RECT 4.395 0.255 4.755 1.075 ;
        RECT 4.975 0.085 5.265 0.905 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor2b_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__nor3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nor3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.740 0.655 2.205 1.665 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.595 1.325 0.880 2.005 ;
        RECT 0.595 0.995 1.075 1.325 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.995 0.425 1.325 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.265 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.647000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 2.280 1.415 2.450 ;
        RECT 0.090 1.495 0.425 2.280 ;
        RECT 1.245 0.825 1.415 2.280 ;
        RECT 0.090 0.655 1.415 0.825 ;
        RECT 0.090 0.385 0.345 0.655 ;
        RECT 1.115 0.385 1.285 0.655 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 1.585 1.835 2.175 2.635 ;
        RECT 0.515 0.085 0.895 0.485 ;
        RECT 1.455 0.085 2.175 0.485 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor3_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__nor3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nor3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.135 1.075 1.015 1.285 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 1.235 1.075 2.275 1.285 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.285 2.935 1.625 ;
        RECT 2.445 1.075 3.310 1.285 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.105 3.990 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.011500 ;
    PORT
      LAYER li1 ;
        RECT 3.180 1.625 3.390 2.125 ;
        RECT 3.180 1.455 3.995 1.625 ;
        RECT 3.480 0.905 3.995 1.455 ;
        RECT 0.535 0.725 3.995 0.905 ;
        RECT 0.535 0.255 0.915 0.725 ;
        RECT 1.475 0.255 1.855 0.725 ;
        RECT 3.050 0.255 3.430 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.150 1.625 0.405 2.465 ;
        RECT 0.625 1.795 0.875 2.635 ;
        RECT 1.095 1.625 1.345 2.465 ;
        RECT 1.565 2.295 3.860 2.465 ;
        RECT 1.565 1.795 1.815 2.295 ;
        RECT 2.035 1.625 2.275 2.125 ;
        RECT 2.710 1.795 2.920 2.295 ;
        RECT 3.610 1.795 3.860 2.295 ;
        RECT 0.150 1.455 2.275 1.625 ;
        RECT 0.090 0.085 0.365 0.905 ;
        RECT 1.135 0.085 1.305 0.555 ;
        RECT 2.075 0.085 2.880 0.555 ;
        RECT 3.650 0.085 3.940 0.555 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor3_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__nor3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nor3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 2.025 1.285 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 3.915 1.445 5.715 1.615 ;
        RECT 3.915 1.285 4.085 1.445 ;
        RECT 2.295 1.075 4.085 1.285 ;
        RECT 5.545 1.285 5.715 1.445 ;
        RECT 5.545 1.075 5.885 1.285 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 4.255 1.075 5.315 1.275 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 6.175 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.828000 ;
    PORT
      LAYER li1 ;
        RECT 3.915 1.965 4.165 2.125 ;
        RECT 4.855 1.965 5.105 2.125 ;
        RECT 3.915 1.955 5.105 1.965 ;
        RECT 3.915 1.785 6.345 1.955 ;
        RECT 6.055 0.905 6.345 1.785 ;
        RECT 0.535 0.725 6.345 0.905 ;
        RECT 0.535 0.255 0.915 0.725 ;
        RECT 1.475 0.255 1.855 0.725 ;
        RECT 2.415 0.255 2.795 0.725 ;
        RECT 3.355 0.255 3.735 0.725 ;
        RECT 4.295 0.255 4.675 0.725 ;
        RECT 5.235 0.255 5.615 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.150 1.625 0.405 2.465 ;
        RECT 0.625 1.795 0.875 2.635 ;
        RECT 1.095 1.625 1.345 2.465 ;
        RECT 1.565 1.795 1.815 2.635 ;
        RECT 2.035 2.085 3.225 2.465 ;
        RECT 2.035 1.625 2.285 2.085 ;
        RECT 0.150 1.455 2.285 1.625 ;
        RECT 2.505 1.625 2.755 1.915 ;
        RECT 2.975 1.795 3.225 2.085 ;
        RECT 3.445 2.295 5.575 2.465 ;
        RECT 3.445 1.625 3.695 2.295 ;
        RECT 4.385 2.135 4.635 2.295 ;
        RECT 5.325 2.135 5.575 2.295 ;
        RECT 5.795 2.125 6.045 2.465 ;
        RECT 2.505 1.455 3.695 1.625 ;
        RECT 0.090 0.085 0.365 0.905 ;
        RECT 1.135 0.085 1.305 0.555 ;
        RECT 2.075 0.085 2.245 0.555 ;
        RECT 3.015 0.085 3.185 0.555 ;
        RECT 3.955 0.085 4.125 0.555 ;
        RECT 4.895 0.085 5.065 0.555 ;
        RECT 5.835 0.085 6.005 0.555 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 2.695 2.125 2.865 2.295 ;
        RECT 5.805 2.125 5.975 2.295 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
      LAYER met1 ;
        RECT 2.635 2.280 2.980 2.335 ;
        RECT 5.695 2.280 6.040 2.335 ;
        RECT 2.635 2.140 6.040 2.280 ;
        RECT 2.635 2.065 2.980 2.140 ;
        RECT 5.695 2.065 6.040 2.140 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor3_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__nor3b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nor3b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.475 0.995 1.815 1.615 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.055 0.995 1.305 1.615 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.985 0.995 2.335 1.615 ;
    END
  END C_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.185 0.335 2.720 1.015 ;
        RECT 0.185 0.105 2.185 0.335 ;
        RECT 0.185 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.759000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.445 0.545 2.455 ;
        RECT 0.085 0.825 0.255 1.445 ;
        RECT 0.085 0.655 1.545 0.825 ;
        RECT 0.085 0.255 0.605 0.655 ;
        RECT 1.375 0.310 1.545 0.655 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 1.715 2.125 2.095 2.635 ;
        RECT 0.715 1.785 2.675 1.955 ;
        RECT 0.715 1.245 0.885 1.785 ;
        RECT 0.425 1.075 0.885 1.245 ;
        RECT 2.505 0.825 2.675 1.785 ;
        RECT 0.775 0.085 1.155 0.485 ;
        RECT 1.715 0.085 2.095 0.825 ;
        RECT 2.380 0.655 2.675 0.825 ;
        RECT 2.380 0.405 2.550 0.655 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor3b_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__nor3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nor3b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.110 1.075 1.015 1.285 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 1.235 1.075 2.200 1.285 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 4.330 1.075 4.915 1.285 ;
    END
  END C_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.335 4.945 1.015 ;
        RECT 0.005 0.105 3.935 0.335 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.979000 ;
    PORT
      LAYER li1 ;
        RECT 2.870 0.905 3.355 2.045 ;
        RECT 0.535 0.725 3.355 0.905 ;
        RECT 0.535 0.255 0.915 0.725 ;
        RECT 1.475 0.255 1.855 0.725 ;
        RECT 2.935 0.255 3.355 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.060 2.805 ;
        RECT 0.090 1.625 0.405 2.465 ;
        RECT 0.625 1.795 0.875 2.635 ;
        RECT 1.095 1.625 1.345 2.465 ;
        RECT 1.565 2.275 3.780 2.465 ;
        RECT 1.565 1.795 1.815 2.275 ;
        RECT 1.995 1.625 2.325 2.035 ;
        RECT 0.090 1.455 2.325 1.625 ;
        RECT 3.535 1.455 3.780 2.275 ;
        RECT 3.990 1.455 4.345 1.870 ;
        RECT 4.565 1.540 4.815 2.635 ;
        RECT 3.990 1.285 4.160 1.455 ;
        RECT 3.535 1.075 4.160 1.285 ;
        RECT 3.990 0.905 4.160 1.075 ;
        RECT 0.090 0.085 0.365 0.905 ;
        RECT 1.135 0.085 1.305 0.555 ;
        RECT 2.075 0.085 2.765 0.555 ;
        RECT 3.575 0.085 3.780 0.895 ;
        RECT 3.990 0.380 4.345 0.905 ;
        RECT 4.565 0.085 4.855 0.825 ;
        RECT 0.000 -0.085 5.060 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor3b_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__nor3b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nor3b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 1.210 1.075 2.770 1.285 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 3.285 1.075 4.700 1.285 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.110 1.075 0.445 1.285 ;
    END
  END C_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 7.165 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.925500 ;
    PORT
      LAYER li1 ;
        RECT 5.375 1.625 5.625 2.125 ;
        RECT 6.315 1.625 6.565 2.125 ;
        RECT 5.375 1.455 7.245 1.625 ;
        RECT 6.905 0.905 7.245 1.455 ;
        RECT 1.005 0.725 7.245 0.905 ;
        RECT 1.005 0.255 1.385 0.725 ;
        RECT 1.945 0.255 2.325 0.725 ;
        RECT 3.405 0.255 3.785 0.725 ;
        RECT 4.345 0.255 4.725 0.725 ;
        RECT 5.285 0.255 5.665 0.725 ;
        RECT 6.225 0.255 6.605 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.360 2.805 ;
        RECT 0.110 1.625 0.405 2.465 ;
        RECT 0.625 1.795 0.875 2.635 ;
        RECT 1.095 1.965 1.345 2.465 ;
        RECT 1.565 2.135 1.815 2.635 ;
        RECT 2.035 1.965 2.285 2.465 ;
        RECT 2.505 2.135 2.755 2.635 ;
        RECT 3.025 2.295 7.035 2.465 ;
        RECT 3.025 2.135 3.275 2.295 ;
        RECT 3.965 2.135 4.215 2.295 ;
        RECT 3.495 1.965 3.745 2.125 ;
        RECT 4.435 1.965 4.685 2.125 ;
        RECT 1.095 1.795 4.685 1.965 ;
        RECT 4.905 1.795 5.155 2.295 ;
        RECT 5.845 1.795 6.095 2.295 ;
        RECT 6.785 1.795 7.035 2.295 ;
        RECT 0.110 1.455 5.155 1.625 ;
        RECT 0.665 0.905 0.835 1.455 ;
        RECT 4.985 1.285 5.155 1.455 ;
        RECT 4.985 1.075 6.720 1.285 ;
        RECT 0.110 0.735 0.835 0.905 ;
        RECT 0.110 0.255 0.445 0.735 ;
        RECT 0.665 0.085 0.835 0.555 ;
        RECT 1.605 0.085 1.775 0.555 ;
        RECT 2.545 0.085 3.235 0.555 ;
        RECT 4.005 0.085 4.175 0.555 ;
        RECT 4.945 0.085 5.115 0.555 ;
        RECT 5.885 0.085 6.055 0.555 ;
        RECT 6.825 0.085 6.995 0.555 ;
        RECT 0.000 -0.085 7.360 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor3b_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__nor4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nor4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.935 0.655 2.205 1.665 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.455 0.995 1.745 2.450 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.965 0.995 1.285 2.450 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.745 0.335 1.325 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.455 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.699000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.665 0.425 2.450 ;
        RECT 0.090 1.495 0.775 1.665 ;
        RECT 0.515 0.825 0.775 1.495 ;
        RECT 0.515 0.655 1.765 0.825 ;
        RECT 0.515 0.385 0.815 0.655 ;
        RECT 1.595 0.385 1.765 0.655 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 2.135 1.835 2.535 2.635 ;
        RECT 0.085 0.085 0.345 0.575 ;
        RECT 1.035 0.085 1.365 0.485 ;
        RECT 2.005 0.085 2.520 0.485 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor4_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__nor4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nor4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.200 1.075 1.015 1.285 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 1.235 1.075 2.140 1.285 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.410 1.075 3.355 1.285 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 3.640 1.075 4.275 1.285 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.855 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.252000 ;
    PORT
      LAYER li1 ;
        RECT 4.040 1.625 4.290 2.125 ;
        RECT 4.040 1.455 4.950 1.625 ;
        RECT 4.615 0.905 4.950 1.455 ;
        RECT 0.570 0.725 4.950 0.905 ;
        RECT 0.570 0.255 0.950 0.725 ;
        RECT 1.510 0.255 1.890 0.725 ;
        RECT 3.010 0.255 3.390 0.725 ;
        RECT 3.950 0.255 4.330 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.060 2.805 ;
        RECT 0.150 1.625 0.405 2.465 ;
        RECT 0.625 1.795 0.875 2.635 ;
        RECT 1.095 1.625 1.345 2.465 ;
        RECT 1.565 2.295 3.315 2.465 ;
        RECT 1.565 1.795 1.815 2.295 ;
        RECT 2.035 1.625 2.285 2.125 ;
        RECT 0.150 1.455 2.285 1.625 ;
        RECT 2.595 1.625 2.845 2.125 ;
        RECT 3.065 1.795 3.315 2.295 ;
        RECT 3.535 2.295 4.725 2.465 ;
        RECT 3.535 1.625 3.785 2.295 ;
        RECT 4.475 1.795 4.725 2.295 ;
        RECT 2.595 1.455 3.785 1.625 ;
        RECT 0.090 0.085 0.365 0.905 ;
        RECT 1.135 0.085 1.305 0.555 ;
        RECT 2.075 0.085 2.805 0.555 ;
        RECT 3.575 0.085 3.745 0.555 ;
        RECT 4.515 0.085 4.805 0.555 ;
        RECT 0.000 -0.085 5.060 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor4_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__nor4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nor4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.740 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.180 1.075 2.025 1.285 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 2.295 1.075 4.470 1.285 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 4.695 1.075 6.305 1.285 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 6.475 1.075 8.045 1.285 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.740 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 8.575 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.930 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.740 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.374000 ;
    PORT
      LAYER li1 ;
        RECT 6.785 1.625 7.035 2.125 ;
        RECT 7.725 1.625 7.975 2.125 ;
        RECT 6.785 1.455 8.630 1.625 ;
        RECT 8.360 0.905 8.630 1.455 ;
        RECT 0.535 0.725 8.630 0.905 ;
        RECT 0.535 0.255 0.915 0.725 ;
        RECT 1.475 0.255 1.855 0.725 ;
        RECT 2.415 0.255 2.795 0.725 ;
        RECT 3.355 0.255 3.735 0.725 ;
        RECT 4.815 0.255 5.195 0.725 ;
        RECT 5.755 0.255 6.135 0.725 ;
        RECT 6.695 0.255 7.075 0.725 ;
        RECT 7.635 0.255 8.015 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.740 2.805 ;
        RECT 0.090 1.625 0.405 2.465 ;
        RECT 0.625 1.795 0.875 2.635 ;
        RECT 1.095 1.625 1.345 2.465 ;
        RECT 1.565 1.795 1.815 2.635 ;
        RECT 2.035 2.295 4.220 2.465 ;
        RECT 2.035 1.625 2.285 2.295 ;
        RECT 0.090 1.455 2.285 1.625 ;
        RECT 2.505 1.625 2.755 2.125 ;
        RECT 2.975 1.795 3.225 2.295 ;
        RECT 3.445 1.625 3.695 2.125 ;
        RECT 3.915 1.795 4.220 2.295 ;
        RECT 4.405 2.295 8.445 2.465 ;
        RECT 4.405 1.795 4.685 2.295 ;
        RECT 4.905 1.625 5.155 2.125 ;
        RECT 5.375 1.795 5.625 2.295 ;
        RECT 5.845 1.625 6.095 2.125 ;
        RECT 6.315 1.795 6.565 2.295 ;
        RECT 7.255 1.795 7.505 2.295 ;
        RECT 8.195 1.795 8.445 2.295 ;
        RECT 2.505 1.455 6.095 1.625 ;
        RECT 0.090 0.085 0.365 0.905 ;
        RECT 1.135 0.085 1.305 0.555 ;
        RECT 2.075 0.085 2.245 0.555 ;
        RECT 3.015 0.085 3.185 0.555 ;
        RECT 3.955 0.085 4.645 0.555 ;
        RECT 5.415 0.085 5.585 0.555 ;
        RECT 6.355 0.085 6.525 0.555 ;
        RECT 7.295 0.085 7.465 0.555 ;
        RECT 8.235 0.085 8.405 0.555 ;
        RECT 0.000 -0.085 8.740 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor4_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__nor4_6
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nor4_6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.420 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.665000 ;
    PORT
      LAYER li1 ;
        RECT 0.505 1.075 2.875 1.285 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.665000 ;
    PORT
      LAYER li1 ;
        RECT 3.325 1.075 5.695 1.285 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.665000 ;
    PORT
      LAYER li1 ;
        RECT 6.665 1.075 9.035 1.285 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.665000 ;
    PORT
      LAYER li1 ;
        RECT 9.395 1.075 11.085 1.285 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 12.420 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 12.365 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 12.610 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 12.420 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.976000 ;
    PORT
      LAYER li1 ;
        RECT 9.605 1.625 9.855 2.125 ;
        RECT 10.545 1.625 10.795 2.125 ;
        RECT 11.445 1.625 11.835 2.125 ;
        RECT 9.605 1.455 11.835 1.625 ;
        RECT 11.445 0.905 11.835 1.455 ;
        RECT 0.585 0.725 11.835 0.905 ;
        RECT 0.585 0.255 0.915 0.725 ;
        RECT 1.525 0.255 1.855 0.725 ;
        RECT 2.465 0.255 2.795 0.725 ;
        RECT 3.405 0.255 3.735 0.725 ;
        RECT 4.345 0.255 4.675 0.725 ;
        RECT 5.285 0.255 5.615 0.725 ;
        RECT 6.745 0.255 7.075 0.725 ;
        RECT 7.685 0.255 8.015 0.725 ;
        RECT 8.625 0.255 8.955 0.725 ;
        RECT 9.565 0.255 9.895 0.725 ;
        RECT 10.505 0.255 10.835 0.725 ;
        RECT 11.445 0.255 11.835 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 12.420 2.805 ;
        RECT 0.115 1.625 0.405 2.465 ;
        RECT 0.625 1.795 0.875 2.635 ;
        RECT 1.095 1.625 1.345 2.465 ;
        RECT 1.565 1.795 1.815 2.635 ;
        RECT 2.035 1.625 2.285 2.465 ;
        RECT 2.505 1.795 2.755 2.635 ;
        RECT 2.975 2.295 6.085 2.465 ;
        RECT 2.975 1.625 3.225 2.295 ;
        RECT 0.115 1.455 3.225 1.625 ;
        RECT 3.445 1.625 3.695 2.125 ;
        RECT 3.915 1.795 4.165 2.295 ;
        RECT 4.385 1.625 4.635 2.125 ;
        RECT 4.855 1.795 5.105 2.295 ;
        RECT 5.325 1.625 5.575 2.125 ;
        RECT 5.795 1.795 6.085 2.295 ;
        RECT 6.275 2.295 12.255 2.465 ;
        RECT 6.275 1.795 6.565 2.295 ;
        RECT 6.785 1.625 7.035 2.125 ;
        RECT 7.255 1.795 7.505 2.295 ;
        RECT 7.725 1.625 7.975 2.125 ;
        RECT 8.195 1.795 8.445 2.295 ;
        RECT 8.665 1.625 8.915 2.125 ;
        RECT 3.445 1.455 8.915 1.625 ;
        RECT 9.135 1.455 9.385 2.295 ;
        RECT 10.075 1.795 10.325 2.295 ;
        RECT 11.015 1.795 11.265 2.295 ;
        RECT 12.005 1.455 12.255 2.295 ;
        RECT 0.115 0.085 0.415 0.905 ;
        RECT 1.085 0.085 1.355 0.555 ;
        RECT 2.025 0.085 2.295 0.555 ;
        RECT 2.965 0.085 3.235 0.555 ;
        RECT 3.905 0.085 4.175 0.555 ;
        RECT 4.845 0.085 5.115 0.555 ;
        RECT 5.785 0.085 6.575 0.555 ;
        RECT 7.245 0.085 7.515 0.555 ;
        RECT 8.185 0.085 8.455 0.555 ;
        RECT 9.125 0.085 9.395 0.555 ;
        RECT 10.065 0.085 10.335 0.555 ;
        RECT 11.005 0.085 11.275 0.555 ;
        RECT 12.005 0.085 12.255 0.905 ;
        RECT 0.000 -0.085 12.420 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor4_6

#--------EOF---------

MACRO sky130_fd_sc_hdll__nor4_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nor4_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.100 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.220000 ;
    PORT
      LAYER li1 ;
        RECT 0.405 1.075 3.795 1.285 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.220000 ;
    PORT
      LAYER li1 ;
        RECT 4.245 1.075 7.635 1.285 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.220000 ;
    PORT
      LAYER li1 ;
        RECT 8.445 1.075 11.835 1.285 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.220000 ;
    PORT
      LAYER li1 ;
        RECT 12.985 1.075 15.355 1.285 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 16.100 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 16.085 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 16.290 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 16.100 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.968000 ;
    PORT
      LAYER li1 ;
        RECT 12.405 1.625 12.655 2.125 ;
        RECT 13.345 1.625 13.595 2.125 ;
        RECT 14.285 1.625 14.535 2.125 ;
        RECT 15.225 1.625 15.475 2.125 ;
        RECT 12.405 1.455 15.475 1.625 ;
        RECT 12.405 0.905 12.815 1.455 ;
        RECT 0.565 0.725 15.515 0.905 ;
        RECT 0.565 0.255 0.895 0.725 ;
        RECT 1.505 0.255 1.835 0.725 ;
        RECT 2.445 0.255 2.775 0.725 ;
        RECT 3.385 0.255 3.715 0.725 ;
        RECT 4.325 0.255 4.655 0.725 ;
        RECT 5.265 0.255 5.595 0.725 ;
        RECT 6.205 0.255 6.535 0.725 ;
        RECT 7.145 0.255 7.475 0.725 ;
        RECT 8.605 0.255 8.935 0.725 ;
        RECT 9.545 0.255 9.875 0.725 ;
        RECT 10.485 0.255 10.815 0.725 ;
        RECT 11.425 0.255 11.755 0.725 ;
        RECT 12.365 0.255 12.695 0.725 ;
        RECT 13.305 0.255 13.635 0.725 ;
        RECT 14.245 0.255 14.575 0.725 ;
        RECT 15.185 0.255 15.515 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 16.100 2.805 ;
        RECT 0.095 1.625 0.425 2.465 ;
        RECT 0.605 1.795 0.855 2.635 ;
        RECT 1.075 1.625 1.325 2.465 ;
        RECT 1.545 1.795 1.795 2.635 ;
        RECT 2.015 1.625 2.265 2.465 ;
        RECT 2.485 1.795 2.735 2.635 ;
        RECT 2.955 1.625 3.205 2.465 ;
        RECT 3.425 1.795 3.675 2.635 ;
        RECT 3.895 2.295 7.945 2.465 ;
        RECT 3.895 1.625 4.145 2.295 ;
        RECT 0.095 1.455 4.145 1.625 ;
        RECT 4.365 1.625 4.615 2.125 ;
        RECT 4.835 1.795 5.085 2.295 ;
        RECT 5.305 1.625 5.555 2.125 ;
        RECT 5.775 1.795 6.025 2.295 ;
        RECT 6.245 1.625 6.495 2.125 ;
        RECT 6.715 1.795 6.965 2.295 ;
        RECT 7.185 1.625 7.435 2.125 ;
        RECT 7.655 1.795 7.945 2.295 ;
        RECT 8.135 2.295 15.995 2.465 ;
        RECT 8.135 1.795 8.425 2.295 ;
        RECT 8.645 1.625 8.895 2.125 ;
        RECT 9.075 1.795 9.365 2.295 ;
        RECT 9.585 1.625 9.835 2.125 ;
        RECT 10.055 1.795 10.305 2.295 ;
        RECT 10.525 1.625 10.775 2.125 ;
        RECT 10.995 1.795 11.245 2.295 ;
        RECT 11.465 1.625 11.715 2.125 ;
        RECT 4.365 1.455 11.715 1.625 ;
        RECT 11.935 1.455 12.185 2.295 ;
        RECT 12.875 1.795 13.125 2.295 ;
        RECT 13.815 1.795 14.065 2.295 ;
        RECT 14.755 1.795 15.005 2.295 ;
        RECT 15.695 1.465 15.995 2.295 ;
        RECT 0.135 0.085 0.395 0.905 ;
        RECT 1.065 0.085 1.335 0.555 ;
        RECT 2.005 0.085 2.275 0.555 ;
        RECT 2.945 0.085 3.215 0.555 ;
        RECT 3.885 0.085 4.155 0.555 ;
        RECT 4.825 0.085 5.095 0.555 ;
        RECT 5.765 0.085 6.035 0.555 ;
        RECT 6.705 0.085 6.975 0.555 ;
        RECT 7.645 0.085 8.435 0.555 ;
        RECT 9.105 0.085 9.375 0.555 ;
        RECT 10.045 0.085 10.315 0.555 ;
        RECT 10.985 0.085 11.255 0.555 ;
        RECT 11.925 0.085 12.195 0.555 ;
        RECT 12.865 0.085 13.135 0.555 ;
        RECT 13.805 0.085 14.075 0.555 ;
        RECT 14.745 0.085 15.015 0.555 ;
        RECT 15.685 0.085 15.965 0.905 ;
        RECT 0.000 -0.085 16.100 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 14.405 2.635 14.575 2.805 ;
        RECT 14.865 2.635 15.035 2.805 ;
        RECT 15.325 2.635 15.495 2.805 ;
        RECT 15.785 2.635 15.955 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
        RECT 14.405 -0.085 14.575 0.085 ;
        RECT 14.865 -0.085 15.035 0.085 ;
        RECT 15.325 -0.085 15.495 0.085 ;
        RECT 15.785 -0.085 15.955 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor4_8

#--------EOF---------

MACRO sky130_fd_sc_hdll__nor4b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nor4b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.175 0.995 2.655 1.615 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.475 0.995 1.935 1.615 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.935 0.995 1.285 1.615 ;
    END
  END C
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 2.825 0.995 3.225 1.615 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.245 0.335 3.430 1.015 ;
        RECT 0.245 0.105 2.865 0.335 ;
        RECT 0.245 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.913500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.825 0.345 2.450 ;
        RECT 0.085 0.655 2.075 0.825 ;
        RECT 0.905 0.300 1.105 0.655 ;
        RECT 1.875 0.310 2.075 0.655 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 2.325 2.185 2.705 2.635 ;
        RECT 0.525 1.795 3.565 2.005 ;
        RECT 0.525 0.995 0.745 1.795 ;
        RECT 3.395 0.825 3.565 1.795 ;
        RECT 0.355 0.085 0.685 0.480 ;
        RECT 1.325 0.085 1.655 0.485 ;
        RECT 2.245 0.085 2.735 0.825 ;
        RECT 3.090 0.655 3.565 0.825 ;
        RECT 3.090 0.405 3.260 0.655 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor4b_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__nor4b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nor4b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.100 1.075 1.340 1.285 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 1.525 1.075 2.650 1.285 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.860 1.075 3.660 1.285 ;
    END
  END C
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 5.615 1.285 5.885 1.955 ;
        RECT 5.205 1.075 5.885 1.285 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.335 5.820 1.015 ;
        RECT 0.005 0.105 4.830 0.335 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.219500 ;
    PORT
      LAYER li1 ;
        RECT 3.980 1.625 4.230 2.125 ;
        RECT 3.980 1.455 4.490 1.625 ;
        RECT 4.065 1.075 4.490 1.455 ;
        RECT 4.065 0.905 4.270 1.075 ;
        RECT 0.515 0.725 4.270 0.905 ;
        RECT 0.515 0.255 0.895 0.725 ;
        RECT 1.455 0.255 1.835 0.725 ;
        RECT 2.950 0.255 3.330 0.725 ;
        RECT 3.890 0.255 4.270 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.085 1.625 0.425 2.465 ;
        RECT 0.645 1.795 0.855 2.635 ;
        RECT 1.075 1.625 1.325 2.465 ;
        RECT 1.545 2.295 3.290 2.465 ;
        RECT 1.545 1.795 1.755 2.295 ;
        RECT 1.925 1.625 2.305 2.125 ;
        RECT 0.085 1.455 2.305 1.625 ;
        RECT 2.475 1.625 2.860 2.125 ;
        RECT 3.080 1.795 3.290 2.295 ;
        RECT 3.510 2.295 4.695 2.465 ;
        RECT 3.510 1.625 3.760 2.295 ;
        RECT 4.450 1.795 4.695 2.295 ;
        RECT 4.865 2.035 5.220 2.450 ;
        RECT 5.440 2.135 5.690 2.635 ;
        RECT 2.475 1.455 3.760 1.625 ;
        RECT 4.865 1.245 5.035 2.035 ;
        RECT 4.720 1.075 5.035 1.245 ;
        RECT 4.865 0.905 5.035 1.075 ;
        RECT 0.085 0.085 0.345 0.905 ;
        RECT 1.115 0.085 1.285 0.555 ;
        RECT 2.055 0.085 2.780 0.555 ;
        RECT 3.550 0.085 3.720 0.555 ;
        RECT 4.490 0.085 4.695 0.895 ;
        RECT 4.865 0.380 5.220 0.905 ;
        RECT 5.440 0.085 5.690 0.825 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor4b_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__nor4b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nor4b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.660 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.395 1.075 2.005 1.285 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 2.275 1.075 4.150 1.285 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 4.385 1.075 6.285 1.285 ;
    END
  END C
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 8.855 1.075 9.550 1.285 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.660 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 9.565 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.850 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.660 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.341500 ;
    PORT
      LAYER li1 ;
        RECT 6.765 1.625 7.015 2.125 ;
        RECT 7.705 1.625 7.955 2.125 ;
        RECT 6.765 1.455 7.955 1.625 ;
        RECT 6.765 0.905 7.250 1.455 ;
        RECT 0.515 0.725 7.995 0.905 ;
        RECT 0.515 0.255 0.895 0.725 ;
        RECT 1.455 0.255 1.835 0.725 ;
        RECT 2.395 0.255 2.775 0.725 ;
        RECT 3.335 0.255 3.715 0.725 ;
        RECT 4.795 0.255 5.175 0.725 ;
        RECT 5.735 0.255 6.115 0.725 ;
        RECT 6.675 0.255 7.055 0.725 ;
        RECT 7.615 0.255 7.995 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.660 2.805 ;
        RECT 0.095 1.625 0.425 2.465 ;
        RECT 0.645 1.795 0.855 2.635 ;
        RECT 1.075 1.625 1.325 2.465 ;
        RECT 1.545 1.795 1.795 2.635 ;
        RECT 2.015 2.295 4.145 2.465 ;
        RECT 2.015 1.625 2.265 2.295 ;
        RECT 0.095 1.455 2.265 1.625 ;
        RECT 2.485 1.625 2.735 2.125 ;
        RECT 2.955 1.795 3.205 2.295 ;
        RECT 3.425 1.625 3.675 2.125 ;
        RECT 3.895 1.795 4.145 2.295 ;
        RECT 4.415 2.295 8.425 2.465 ;
        RECT 4.415 1.795 4.665 2.295 ;
        RECT 4.885 1.625 5.135 2.125 ;
        RECT 5.355 1.795 5.605 2.295 ;
        RECT 5.825 1.625 6.075 2.125 ;
        RECT 2.485 1.455 6.075 1.625 ;
        RECT 6.295 1.455 6.545 2.295 ;
        RECT 7.235 1.795 7.485 2.295 ;
        RECT 8.175 1.795 8.425 2.295 ;
        RECT 8.650 1.625 8.985 2.465 ;
        RECT 8.270 1.455 8.985 1.625 ;
        RECT 9.205 1.455 9.435 2.635 ;
        RECT 8.270 1.285 8.440 1.455 ;
        RECT 7.420 1.075 8.440 1.285 ;
        RECT 8.270 0.905 8.440 1.075 ;
        RECT 0.175 0.085 0.345 0.895 ;
        RECT 8.270 0.735 8.985 0.905 ;
        RECT 1.115 0.085 1.285 0.555 ;
        RECT 2.055 0.085 2.225 0.555 ;
        RECT 2.995 0.085 3.165 0.555 ;
        RECT 3.935 0.085 4.625 0.555 ;
        RECT 5.395 0.085 5.565 0.555 ;
        RECT 6.335 0.085 6.505 0.555 ;
        RECT 7.275 0.085 7.445 0.555 ;
        RECT 8.215 0.085 8.385 0.555 ;
        RECT 8.610 0.255 8.985 0.735 ;
        RECT 9.205 0.085 9.435 0.905 ;
        RECT 0.000 -0.085 9.660 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor4b_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__nor4bb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nor4bb_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 3.360 0.995 3.665 1.705 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.820 0.995 3.130 2.410 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.430 0.995 0.830 1.695 ;
    END
  END C_N
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.000 0.995 1.340 1.325 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.045 0.335 3.980 1.015 ;
        RECT 0.150 -0.085 0.320 0.335 ;
        RECT 1.530 0.105 3.980 0.335 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.660000 ;
    PORT
      LAYER li1 ;
        RECT 1.575 1.955 2.210 2.125 ;
        RECT 1.960 0.825 2.210 1.955 ;
        RECT 1.960 0.655 3.340 0.825 ;
        RECT 2.170 0.300 2.370 0.655 ;
        RECT 3.140 0.310 3.340 0.655 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.085 2.070 0.345 2.455 ;
        RECT 0.515 2.240 0.895 2.635 ;
        RECT 1.135 2.295 2.615 2.465 ;
        RECT 1.135 2.070 1.305 2.295 ;
        RECT 0.085 1.885 1.305 2.070 ;
        RECT 0.085 0.825 0.260 1.885 ;
        RECT 1.100 1.525 1.790 1.715 ;
        RECT 1.620 0.825 1.790 1.525 ;
        RECT 2.380 0.995 2.615 2.295 ;
        RECT 3.510 1.875 3.990 2.635 ;
        RECT 0.085 0.450 0.405 0.825 ;
        RECT 0.705 0.085 0.875 0.825 ;
        RECT 1.175 0.655 1.790 0.825 ;
        RECT 1.175 0.450 1.345 0.655 ;
        RECT 1.620 0.085 1.950 0.480 ;
        RECT 2.590 0.085 2.920 0.485 ;
        RECT 3.510 0.085 3.990 0.825 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor4bb_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__nor4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nor4bb_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 5.465 1.075 6.330 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 4.400 1.075 5.295 1.275 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.000 0.995 1.270 1.325 ;
    END
  END C_N
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.995 0.830 1.695 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.335 6.410 1.015 ;
        RECT 0.145 -0.085 0.315 0.335 ;
        RECT 1.505 0.105 6.410 0.335 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.219500 ;
    PORT
      LAYER li1 ;
        RECT 3.035 1.445 4.230 1.705 ;
        RECT 3.810 0.905 4.230 1.445 ;
        RECT 2.095 0.725 5.835 0.905 ;
        RECT 2.095 0.255 2.475 0.725 ;
        RECT 3.035 0.255 3.415 0.725 ;
        RECT 4.515 0.255 4.895 0.725 ;
        RECT 5.455 0.255 5.835 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.085 2.055 0.345 2.455 ;
        RECT 0.515 2.240 0.895 2.635 ;
        RECT 1.675 2.225 3.885 2.465 ;
        RECT 4.095 2.215 5.325 2.465 ;
        RECT 0.085 1.885 1.950 2.055 ;
        RECT 0.085 0.825 0.255 1.885 ;
        RECT 1.045 1.525 1.610 1.715 ;
        RECT 1.440 1.245 1.610 1.525 ;
        RECT 1.780 1.585 1.950 1.885 ;
        RECT 2.145 1.875 4.895 2.045 ;
        RECT 1.780 1.415 2.865 1.585 ;
        RECT 4.605 1.455 4.895 1.875 ;
        RECT 5.115 1.625 5.325 2.215 ;
        RECT 5.545 1.795 5.755 2.635 ;
        RECT 5.925 1.625 6.305 2.465 ;
        RECT 5.115 1.455 6.305 1.625 ;
        RECT 2.695 1.275 2.865 1.415 ;
        RECT 1.440 1.075 2.475 1.245 ;
        RECT 2.695 1.075 3.640 1.275 ;
        RECT 1.440 0.825 1.610 1.075 ;
        RECT 0.085 0.450 0.465 0.825 ;
        RECT 0.685 0.085 0.855 0.825 ;
        RECT 1.155 0.655 1.610 0.825 ;
        RECT 1.155 0.450 1.350 0.655 ;
        RECT 1.595 0.085 1.925 0.480 ;
        RECT 2.695 0.085 2.865 0.555 ;
        RECT 3.635 0.085 4.345 0.555 ;
        RECT 5.115 0.085 5.285 0.555 ;
        RECT 6.055 0.085 6.330 0.905 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor4bb_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__nor4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nor4bb_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.120 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 8.075 1.075 10.010 1.285 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 5.650 1.075 7.805 1.285 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.110 1.075 0.445 1.365 ;
    END
  END C_N
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.075 1.395 1.325 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.120 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.105 10.095 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.310 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.120 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.374000 ;
    PORT
      LAYER li1 ;
        RECT 1.940 1.415 3.435 1.705 ;
        RECT 3.265 0.905 3.435 1.415 ;
        RECT 2.035 0.725 9.515 0.905 ;
        RECT 2.035 0.255 2.415 0.725 ;
        RECT 2.975 0.255 3.355 0.725 ;
        RECT 3.915 0.255 4.295 0.725 ;
        RECT 4.855 0.255 5.235 0.725 ;
        RECT 6.315 0.255 6.695 0.725 ;
        RECT 7.255 0.255 7.635 0.725 ;
        RECT 8.195 0.255 8.575 0.725 ;
        RECT 9.135 0.255 9.515 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.120 2.805 ;
        RECT 0.085 2.045 0.365 2.465 ;
        RECT 0.535 2.215 0.915 2.635 ;
        RECT 1.615 2.295 5.695 2.465 ;
        RECT 1.615 2.215 3.825 2.295 ;
        RECT 0.085 1.875 3.825 2.045 ;
        RECT 0.085 1.535 0.835 1.875 ;
        RECT 1.005 1.535 1.735 1.705 ;
        RECT 0.665 0.895 0.835 1.535 ;
        RECT 1.565 1.245 1.735 1.535 ;
        RECT 3.655 1.285 3.825 1.875 ;
        RECT 4.045 1.625 4.255 2.125 ;
        RECT 4.475 1.795 4.725 2.295 ;
        RECT 4.945 1.625 5.195 2.125 ;
        RECT 5.415 1.795 5.695 2.295 ;
        RECT 5.880 2.295 8.065 2.465 ;
        RECT 5.880 1.795 6.185 2.295 ;
        RECT 6.405 1.625 6.655 2.125 ;
        RECT 6.875 1.795 7.125 2.295 ;
        RECT 7.345 1.625 7.595 2.125 ;
        RECT 4.045 1.455 7.595 1.625 ;
        RECT 7.815 1.625 8.065 2.295 ;
        RECT 8.285 1.795 8.535 2.635 ;
        RECT 8.755 1.625 9.005 2.465 ;
        RECT 9.225 1.795 9.475 2.635 ;
        RECT 9.695 1.625 10.010 2.465 ;
        RECT 7.815 1.455 10.010 1.625 ;
        RECT 1.565 1.075 3.095 1.245 ;
        RECT 3.655 1.075 5.405 1.285 ;
        RECT 1.565 0.905 1.735 1.075 ;
        RECT 0.085 0.725 0.835 0.895 ;
        RECT 1.005 0.735 1.735 0.905 ;
        RECT 0.085 0.255 0.445 0.725 ;
        RECT 0.665 0.085 0.835 0.555 ;
        RECT 1.005 0.255 1.385 0.735 ;
        RECT 1.695 0.085 1.865 0.555 ;
        RECT 2.635 0.085 2.805 0.555 ;
        RECT 3.575 0.085 3.745 0.555 ;
        RECT 4.515 0.085 4.685 0.555 ;
        RECT 5.455 0.085 6.145 0.555 ;
        RECT 6.915 0.085 7.085 0.555 ;
        RECT 7.855 0.085 8.025 0.555 ;
        RECT 8.795 0.085 8.965 0.555 ;
        RECT 9.735 0.085 10.010 0.905 ;
        RECT 0.000 -0.085 10.120 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor4bb_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__o2bb2a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o2bb2a_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.820 1.075 1.320 1.275 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.490 0.905 1.715 1.100 ;
        RECT 1.015 0.735 1.715 0.905 ;
        RECT 1.015 0.380 1.300 0.735 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 3.705 1.075 4.055 1.645 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 3.335 1.325 3.535 2.425 ;
        RECT 2.720 1.075 3.535 1.325 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.785 0.980 1.015 ;
        RECT 0.005 0.105 4.135 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.471500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.795 0.345 2.465 ;
        RECT 0.085 0.825 0.260 1.795 ;
        RECT 0.085 0.255 0.425 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.515 2.235 0.895 2.635 ;
        RECT 1.865 2.235 2.265 2.635 ;
        RECT 2.555 2.055 2.935 2.290 ;
        RECT 0.705 1.885 2.935 2.055 ;
        RECT 0.705 1.615 0.875 1.885 ;
        RECT 0.430 1.445 0.875 1.615 ;
        RECT 1.045 1.495 2.160 1.715 ;
        RECT 0.430 0.995 0.650 1.445 ;
        RECT 1.885 1.355 2.160 1.495 ;
        RECT 2.330 1.495 2.935 1.885 ;
        RECT 3.705 1.815 4.055 2.635 ;
        RECT 0.670 0.085 0.840 0.750 ;
        RECT 1.885 0.565 2.055 1.355 ;
        RECT 2.330 1.245 2.500 1.495 ;
        RECT 2.305 1.075 2.500 1.245 ;
        RECT 2.305 0.690 2.475 1.075 ;
        RECT 1.560 0.395 2.055 0.565 ;
        RECT 2.225 0.320 2.475 0.690 ;
        RECT 2.695 0.725 4.055 0.905 ;
        RECT 2.695 0.320 2.945 0.725 ;
        RECT 3.135 0.085 3.485 0.555 ;
        RECT 3.665 0.320 4.055 0.725 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o2bb2a_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__o2bb2a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o2bb2a_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 1.315 1.075 1.835 1.275 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 2.005 0.905 2.225 1.100 ;
        RECT 1.520 0.735 2.225 0.905 ;
        RECT 1.520 0.380 1.885 0.735 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 4.000 1.075 4.465 1.645 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 3.655 1.915 3.995 2.425 ;
        RECT 3.655 1.325 3.825 1.915 ;
        RECT 3.220 1.075 3.825 1.325 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.785 1.460 1.015 ;
        RECT 0.005 0.105 4.495 0.785 ;
        RECT 0.135 -0.085 0.305 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.498000 ;
    PORT
      LAYER li1 ;
        RECT 0.535 1.795 0.840 2.465 ;
        RECT 0.535 0.825 0.755 1.795 ;
        RECT 0.535 0.255 0.920 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.110 1.410 0.365 2.635 ;
        RECT 1.010 2.235 1.390 2.635 ;
        RECT 2.360 2.235 2.765 2.635 ;
        RECT 3.035 2.055 3.435 2.425 ;
        RECT 1.200 1.885 3.435 2.055 ;
        RECT 1.200 1.615 1.370 1.885 ;
        RECT 0.925 1.445 1.370 1.615 ;
        RECT 1.540 1.495 2.660 1.715 ;
        RECT 0.925 0.995 1.145 1.445 ;
        RECT 2.395 1.355 2.660 1.495 ;
        RECT 2.830 1.495 3.435 1.885 ;
        RECT 4.165 1.815 4.480 2.635 ;
        RECT 0.110 0.085 0.365 0.910 ;
        RECT 1.135 0.085 1.305 0.750 ;
        RECT 2.395 0.565 2.565 1.355 ;
        RECT 2.830 1.245 3.000 1.495 ;
        RECT 2.810 1.075 3.000 1.245 ;
        RECT 2.810 0.690 2.980 1.075 ;
        RECT 2.055 0.395 2.565 0.565 ;
        RECT 2.735 0.320 2.980 0.690 ;
        RECT 3.205 0.725 4.405 0.905 ;
        RECT 3.205 0.320 3.435 0.725 ;
        RECT 3.675 0.085 3.845 0.555 ;
        RECT 4.015 0.320 4.405 0.725 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o2bb2a_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__o2bb2a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o2bb2a_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.820 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 3.615 1.445 5.465 1.615 ;
        RECT 3.615 1.075 3.995 1.445 ;
        RECT 5.055 1.075 5.465 1.445 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 4.165 1.075 4.885 1.275 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.445 2.095 1.615 ;
        RECT 0.085 1.075 0.625 1.445 ;
        RECT 1.715 1.075 2.095 1.445 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.855 1.075 1.445 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.820 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 7.615 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.010 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.820 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.028500 ;
    PORT
      LAYER li1 ;
        RECT 5.825 1.955 6.075 2.465 ;
        RECT 6.765 1.955 7.015 2.465 ;
        RECT 5.825 1.785 7.015 1.955 ;
        RECT 6.765 1.655 7.015 1.785 ;
        RECT 6.765 1.415 7.710 1.655 ;
        RECT 7.405 0.905 7.710 1.415 ;
        RECT 5.735 0.725 7.710 0.905 ;
        RECT 5.735 0.275 6.115 0.725 ;
        RECT 6.675 0.275 7.055 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.820 2.805 ;
        RECT 0.140 1.795 0.345 2.635 ;
        RECT 0.605 2.295 1.795 2.465 ;
        RECT 0.605 1.785 0.855 2.295 ;
        RECT 1.545 2.125 1.795 2.295 ;
        RECT 2.015 2.125 2.265 2.635 ;
        RECT 1.075 1.955 1.325 2.125 ;
        RECT 2.485 1.965 2.775 2.465 ;
        RECT 2.995 2.135 3.725 2.635 ;
        RECT 4.415 2.135 4.665 2.635 ;
        RECT 3.945 1.965 4.195 2.125 ;
        RECT 4.885 1.965 5.135 2.465 ;
        RECT 2.485 1.955 2.865 1.965 ;
        RECT 1.075 1.785 2.865 1.955 ;
        RECT 2.265 1.415 2.865 1.785 ;
        RECT 3.255 1.785 5.135 1.965 ;
        RECT 5.355 1.795 5.605 2.635 ;
        RECT 6.295 2.165 6.545 2.635 ;
        RECT 7.235 1.825 7.485 2.635 ;
        RECT 2.265 1.075 2.695 1.415 ;
        RECT 3.255 1.245 3.445 1.785 ;
        RECT 2.865 1.075 3.445 1.245 ;
        RECT 5.665 1.245 6.005 1.615 ;
        RECT 5.665 1.075 7.085 1.245 ;
        RECT 0.095 0.735 2.225 0.905 ;
        RECT 0.095 0.725 1.365 0.735 ;
        RECT 0.095 0.255 0.425 0.725 ;
        RECT 0.645 0.085 0.815 0.555 ;
        RECT 0.985 0.255 1.365 0.725 ;
        RECT 1.585 0.085 1.755 0.555 ;
        RECT 1.925 0.475 2.225 0.735 ;
        RECT 2.395 0.815 2.695 1.075 ;
        RECT 3.255 0.905 3.445 1.075 ;
        RECT 2.395 0.645 2.775 0.815 ;
        RECT 3.255 0.725 4.705 0.905 ;
        RECT 4.325 0.645 4.705 0.725 ;
        RECT 1.925 0.255 3.245 0.475 ;
        RECT 3.515 0.085 3.685 0.555 ;
        RECT 4.925 0.475 5.175 0.895 ;
        RECT 3.855 0.305 5.175 0.475 ;
        RECT 5.395 0.085 5.565 0.895 ;
        RECT 6.335 0.085 6.505 0.555 ;
        RECT 7.275 0.085 7.445 0.555 ;
        RECT 0.000 -0.085 7.820 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 2.695 1.435 2.865 1.605 ;
        RECT 5.725 1.445 5.895 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
      LAYER met1 ;
        RECT 2.635 1.600 2.975 1.635 ;
        RECT 5.665 1.600 5.960 1.645 ;
        RECT 2.635 1.460 5.960 1.600 ;
        RECT 2.635 1.385 2.975 1.460 ;
        RECT 5.665 1.395 5.960 1.460 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o2bb2a_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__o2bb2ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o2bb2ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.435 1.285 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.995 1.100 1.325 ;
        RECT 0.605 0.280 0.825 0.995 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.865 1.075 3.245 1.285 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.275 2.615 2.425 ;
        RECT 2.150 1.075 2.615 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.330 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.485500 ;
    PORT
      LAYER li1 ;
        RECT 1.950 1.665 2.275 2.465 ;
        RECT 1.760 1.445 2.275 1.665 ;
        RECT 1.760 0.790 1.930 1.445 ;
        RECT 1.610 0.430 1.930 0.790 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.150 1.455 0.400 2.635 ;
        RECT 0.620 1.665 0.870 2.465 ;
        RECT 1.090 1.835 1.780 2.635 ;
        RECT 0.620 1.495 1.440 1.665 ;
        RECT 1.270 1.325 1.440 1.495 ;
        RECT 2.950 1.455 3.200 2.635 ;
        RECT 1.270 0.995 1.580 1.325 ;
        RECT 1.270 0.825 1.440 0.995 ;
        RECT 0.090 0.085 0.425 0.815 ;
        RECT 1.000 0.280 1.440 0.825 ;
        RECT 2.100 0.725 3.240 0.905 ;
        RECT 2.100 0.425 2.350 0.725 ;
        RECT 2.520 0.085 2.690 0.555 ;
        RECT 2.860 0.275 3.240 0.725 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o2bb2ai_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__o2bb2ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o2bb2ai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.445 2.145 1.615 ;
        RECT 0.090 1.075 0.675 1.445 ;
        RECT 1.765 1.075 2.145 1.445 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.845 1.075 1.500 1.275 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 3.650 1.445 5.460 1.615 ;
        RECT 3.650 1.075 4.040 1.445 ;
        RECT 5.130 1.075 5.460 1.445 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 4.260 1.075 4.900 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.750 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.788000 ;
    PORT
      LAYER li1 ;
        RECT 2.895 1.955 3.235 2.465 ;
        RECT 4.430 1.955 4.680 2.125 ;
        RECT 2.895 1.785 4.680 1.955 ;
        RECT 2.895 1.075 3.465 1.785 ;
        RECT 2.895 0.645 3.275 1.075 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.150 1.795 0.400 2.635 ;
        RECT 0.625 1.965 0.875 2.465 ;
        RECT 1.095 2.135 1.345 2.635 ;
        RECT 2.035 2.135 2.725 2.635 ;
        RECT 3.455 2.125 3.740 2.635 ;
        RECT 3.960 2.295 5.150 2.465 ;
        RECT 3.960 2.125 4.210 2.295 ;
        RECT 0.625 1.785 2.485 1.965 ;
        RECT 4.900 1.785 5.150 2.295 ;
        RECT 5.415 1.795 5.620 2.635 ;
        RECT 2.315 1.325 2.485 1.785 ;
        RECT 2.315 0.995 2.725 1.325 ;
        RECT 2.315 0.905 2.485 0.995 ;
        RECT 0.195 0.085 0.365 0.895 ;
        RECT 0.535 0.475 0.835 0.895 ;
        RECT 1.005 0.725 2.485 0.905 ;
        RECT 3.495 0.735 5.660 0.905 ;
        RECT 1.005 0.645 1.385 0.725 ;
        RECT 0.535 0.305 1.855 0.475 ;
        RECT 2.035 0.085 2.205 0.555 ;
        RECT 2.475 0.475 2.725 0.555 ;
        RECT 3.495 0.475 3.780 0.735 ;
        RECT 4.340 0.725 5.660 0.735 ;
        RECT 2.475 0.255 3.780 0.475 ;
        RECT 4.000 0.085 4.170 0.555 ;
        RECT 4.340 0.255 4.720 0.725 ;
        RECT 4.940 0.085 5.110 0.555 ;
        RECT 5.280 0.255 5.660 0.725 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o2bb2ai_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__o2bb2ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o2bb2ai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.040 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 2.295 1.075 3.905 1.285 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.075 2.025 1.285 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 8.845 1.075 10.940 1.285 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 7.065 1.075 8.675 1.285 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.040 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 10.945 1.015 ;
        RECT 0.135 -0.085 0.305 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 11.230 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.040 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.608500 ;
    PORT
      LAYER li1 ;
        RECT 4.875 1.625 5.125 2.465 ;
        RECT 5.815 1.625 6.065 2.465 ;
        RECT 7.275 1.625 7.525 2.125 ;
        RECT 8.215 1.625 8.465 2.125 ;
        RECT 4.875 1.455 8.465 1.625 ;
        RECT 6.475 0.905 6.805 1.455 ;
        RECT 4.865 0.645 6.805 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 11.040 2.805 ;
        RECT 0.155 1.795 0.405 2.635 ;
        RECT 0.625 1.625 0.875 2.465 ;
        RECT 1.095 1.795 1.345 2.635 ;
        RECT 1.565 1.625 1.815 2.465 ;
        RECT 2.035 1.795 2.285 2.635 ;
        RECT 2.505 1.625 2.755 2.465 ;
        RECT 2.975 1.795 3.225 2.635 ;
        RECT 3.445 1.625 3.695 2.465 ;
        RECT 3.915 1.795 4.655 2.635 ;
        RECT 5.345 1.795 5.595 2.635 ;
        RECT 6.285 1.795 6.535 2.635 ;
        RECT 6.775 2.295 8.935 2.465 ;
        RECT 6.775 1.795 7.055 2.295 ;
        RECT 7.745 1.795 7.995 2.295 ;
        RECT 8.685 1.625 8.935 2.295 ;
        RECT 9.155 1.795 9.405 2.635 ;
        RECT 9.625 1.625 9.875 2.465 ;
        RECT 10.095 1.795 10.345 2.635 ;
        RECT 10.565 1.625 10.875 2.465 ;
        RECT 0.085 1.455 4.315 1.625 ;
        RECT 8.685 1.455 10.875 1.625 ;
        RECT 0.085 0.905 0.255 1.455 ;
        RECT 4.145 1.285 4.315 1.455 ;
        RECT 4.145 1.075 6.305 1.285 ;
        RECT 0.085 0.645 1.855 0.905 ;
        RECT 2.075 0.725 4.205 0.905 ;
        RECT 2.075 0.475 2.325 0.725 ;
        RECT 0.100 0.255 2.325 0.475 ;
        RECT 2.545 0.085 2.715 0.555 ;
        RECT 2.885 0.255 3.265 0.725 ;
        RECT 3.485 0.085 3.655 0.555 ;
        RECT 3.825 0.255 4.205 0.725 ;
        RECT 4.460 0.475 4.645 0.835 ;
        RECT 6.975 0.735 10.855 0.905 ;
        RECT 6.975 0.475 7.145 0.735 ;
        RECT 7.655 0.725 10.855 0.735 ;
        RECT 4.460 0.255 7.145 0.475 ;
        RECT 7.315 0.085 7.485 0.555 ;
        RECT 7.655 0.255 8.035 0.725 ;
        RECT 8.255 0.085 8.425 0.555 ;
        RECT 8.595 0.255 8.975 0.725 ;
        RECT 9.195 0.085 9.365 0.555 ;
        RECT 9.535 0.255 9.915 0.725 ;
        RECT 10.135 0.085 10.305 0.555 ;
        RECT 10.475 0.255 10.855 0.725 ;
        RECT 0.000 -0.085 11.040 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o2bb2ai_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__o21a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o21a_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.325 1.075 2.675 1.615 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.985 1.275 2.155 2.390 ;
        RECT 1.725 1.075 2.155 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.055 1.075 1.555 1.305 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.800 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.472000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.030 0.365 2.465 ;
        RECT 0.085 0.255 0.425 1.030 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.535 1.860 1.265 2.635 ;
        RECT 1.480 1.690 1.810 2.465 ;
        RECT 2.380 1.915 3.100 2.635 ;
        RECT 0.600 1.475 1.810 1.690 ;
        RECT 0.600 0.905 0.885 1.475 ;
        RECT 0.600 0.715 1.385 0.905 ;
        RECT 0.615 0.085 0.785 0.545 ;
        RECT 1.025 0.255 1.385 0.715 ;
        RECT 1.555 0.715 2.710 0.905 ;
        RECT 1.555 0.555 1.765 0.715 ;
        RECT 1.980 0.085 2.150 0.545 ;
        RECT 2.380 0.255 2.710 0.715 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o21a_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__o21a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o21a_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 3.275 0.995 3.535 1.450 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.800 1.400 3.075 1.985 ;
        RECT 2.320 1.025 3.075 1.400 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.525 1.010 1.955 1.615 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.625 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.506250 ;
    PORT
      LAYER li1 ;
        RECT 0.530 0.255 0.825 2.465 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.090 1.635 0.345 2.635 ;
        RECT 0.995 2.185 1.895 2.635 ;
        RECT 2.115 2.005 2.375 2.465 ;
        RECT 1.185 1.785 2.375 2.005 ;
        RECT 1.185 1.330 1.355 1.785 ;
        RECT 3.245 1.650 3.530 2.635 ;
        RECT 0.105 0.085 0.345 0.885 ;
        RECT 0.995 0.840 1.355 1.330 ;
        RECT 0.995 0.635 1.895 0.840 ;
        RECT 0.995 0.085 1.375 0.465 ;
        RECT 1.565 0.255 1.895 0.635 ;
        RECT 2.115 0.635 3.530 0.825 ;
        RECT 2.115 0.465 2.325 0.635 ;
        RECT 3.255 0.495 3.530 0.635 ;
        RECT 2.495 0.085 3.035 0.465 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o21a_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__o21a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o21a_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 3.760 1.495 5.880 1.705 ;
        RECT 3.760 0.990 4.115 1.495 ;
        RECT 5.410 0.995 5.880 1.495 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 4.420 0.995 5.070 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.735 1.075 3.485 1.615 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.925 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.029000 ;
    PORT
      LAYER li1 ;
        RECT 1.015 1.700 1.205 2.465 ;
        RECT 1.975 1.700 2.155 2.465 ;
        RECT 0.090 1.530 2.155 1.700 ;
        RECT 0.090 0.805 0.350 1.530 ;
        RECT 0.090 0.635 1.865 0.805 ;
        RECT 0.645 0.615 1.865 0.635 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.415 1.870 0.795 2.635 ;
        RECT 1.375 1.870 1.755 2.635 ;
        RECT 2.335 2.255 2.735 2.635 ;
        RECT 2.955 2.105 3.195 2.465 ;
        RECT 3.515 2.275 3.845 2.635 ;
        RECT 4.495 2.105 4.875 2.445 ;
        RECT 2.955 2.085 4.875 2.105 ;
        RECT 2.325 1.875 4.875 2.085 ;
        RECT 5.455 1.935 5.865 2.635 ;
        RECT 2.325 1.830 3.195 1.875 ;
        RECT 2.325 1.335 2.565 1.830 ;
        RECT 0.520 0.995 2.565 1.335 ;
        RECT 2.315 0.870 2.565 0.995 ;
        RECT 2.315 0.655 3.385 0.870 ;
        RECT 3.555 0.615 5.835 0.785 ;
        RECT 3.555 0.485 3.885 0.615 ;
        RECT 0.095 0.085 0.425 0.465 ;
        RECT 1.055 0.085 1.385 0.445 ;
        RECT 2.015 0.085 2.345 0.465 ;
        RECT 2.585 0.255 3.885 0.485 ;
        RECT 4.055 0.085 4.395 0.445 ;
        RECT 4.975 0.085 5.355 0.445 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o21a_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__o21ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o21ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.995 0.410 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.580 1.325 0.835 2.375 ;
        RECT 0.580 0.995 1.075 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.223500 ;
    PORT
      LAYER li1 ;
        RECT 1.655 1.295 2.215 1.655 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.270 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.752250 ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.505 1.415 2.465 ;
        RECT 1.245 1.125 1.415 1.505 ;
        RECT 1.245 0.955 2.110 1.125 ;
        RECT 1.645 0.275 2.110 0.955 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.090 1.495 0.410 2.635 ;
        RECT 1.645 1.835 2.110 2.635 ;
        RECT 0.090 0.615 1.405 0.785 ;
        RECT 0.090 0.265 0.380 0.615 ;
        RECT 0.625 0.085 1.005 0.445 ;
        RECT 1.175 0.310 1.405 0.615 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o21ai_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__o21ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o21ai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.120 1.445 2.295 1.615 ;
        RECT 0.120 1.055 0.450 1.445 ;
        RECT 1.750 1.075 2.295 1.445 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.670 1.075 1.570 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 3.280 0.765 3.570 1.400 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.015 0.105 3.620 1.015 ;
        RECT 0.140 -0.085 0.310 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.814500 ;
    PORT
      LAYER li1 ;
        RECT 1.095 1.965 1.395 2.125 ;
        RECT 2.695 1.965 3.110 2.465 ;
        RECT 1.095 1.785 3.110 1.965 ;
        RECT 2.695 0.595 3.110 1.785 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.105 1.785 0.435 2.635 ;
        RECT 0.655 2.295 1.865 2.465 ;
        RECT 0.655 1.785 0.875 2.295 ;
        RECT 1.675 2.135 1.865 2.295 ;
        RECT 2.060 2.175 2.440 2.635 ;
        RECT 3.280 1.570 3.530 2.635 ;
        RECT 0.105 0.715 2.465 0.885 ;
        RECT 0.105 0.255 0.435 0.715 ;
        RECT 0.665 0.085 0.835 0.545 ;
        RECT 1.015 0.255 1.395 0.715 ;
        RECT 1.675 0.085 1.845 0.545 ;
        RECT 2.135 0.425 2.465 0.715 ;
        RECT 3.280 0.425 3.530 0.595 ;
        RECT 2.135 0.255 3.530 0.425 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o21ai_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__o21ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o21ai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.625 1.515 4.095 1.685 ;
        RECT 0.625 1.320 1.625 1.515 ;
        RECT 0.125 1.015 1.625 1.320 ;
        RECT 3.795 0.990 4.095 1.515 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 2.185 1.070 3.625 1.345 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 4.305 1.015 5.600 1.275 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.030 0.105 6.360 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.661500 ;
    PORT
      LAYER li1 ;
        RECT 4.530 2.085 4.740 2.465 ;
        RECT 5.510 2.085 5.700 2.465 ;
        RECT 4.530 2.025 5.700 2.085 ;
        RECT 1.990 1.855 5.700 2.025 ;
        RECT 4.335 1.700 5.700 1.855 ;
        RECT 4.335 1.445 6.330 1.700 ;
        RECT 5.920 0.845 6.330 1.445 ;
        RECT 4.430 0.615 6.330 0.845 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.120 1.820 0.405 2.635 ;
        RECT 0.625 2.085 0.860 2.465 ;
        RECT 1.030 2.255 1.410 2.635 ;
        RECT 1.630 2.275 3.810 2.465 ;
        RECT 1.630 2.085 1.820 2.275 ;
        RECT 4.030 2.195 4.310 2.635 ;
        RECT 4.910 2.255 5.290 2.635 ;
        RECT 0.625 1.915 1.820 2.085 ;
        RECT 5.870 1.880 6.250 2.635 ;
        RECT 0.120 0.615 4.260 0.820 ;
        RECT 4.030 0.445 4.260 0.615 ;
        RECT 0.550 0.085 0.930 0.445 ;
        RECT 1.510 0.085 1.890 0.445 ;
        RECT 2.470 0.085 2.850 0.445 ;
        RECT 3.430 0.085 3.810 0.445 ;
        RECT 4.030 0.255 6.250 0.445 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o21ai_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__o21ba_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o21ba_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 3.020 1.075 3.570 1.285 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.230 1.075 2.850 1.285 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.030 0.995 1.380 1.325 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.085 0.105 3.660 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.480 0.425 2.465 ;
        RECT 0.085 0.825 0.340 1.480 ;
        RECT 0.085 0.450 0.445 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.595 2.205 1.005 2.635 ;
        RECT 1.770 2.215 2.100 2.635 ;
        RECT 2.280 2.035 2.585 2.465 ;
        RECT 0.645 1.865 2.585 2.035 ;
        RECT 0.645 1.325 0.860 1.865 ;
        RECT 1.075 1.525 1.720 1.695 ;
        RECT 0.510 0.995 0.860 1.325 ;
        RECT 1.550 0.825 1.720 1.525 ;
        RECT 0.675 0.085 0.845 0.825 ;
        RECT 1.210 0.655 1.720 0.825 ;
        RECT 1.890 1.455 2.585 1.865 ;
        RECT 3.170 1.535 3.550 2.635 ;
        RECT 1.210 0.450 1.380 0.655 ;
        RECT 1.890 0.255 2.060 1.455 ;
        RECT 2.280 0.735 3.565 0.905 ;
        RECT 2.280 0.255 2.610 0.735 ;
        RECT 2.830 0.085 3.000 0.555 ;
        RECT 3.235 0.270 3.565 0.735 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o21ba_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__o21ba_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o21ba_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 3.350 1.075 3.895 1.625 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.645 1.075 3.180 1.285 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.325 0.825 1.695 ;
        RECT 0.425 0.995 0.825 1.325 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.335 3.975 1.015 ;
        RECT 0.145 0.105 3.975 0.335 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.571750 ;
    PORT
      LAYER li1 ;
        RECT 0.995 1.495 1.455 1.695 ;
        RECT 0.995 0.465 1.235 1.495 ;
        RECT 0.995 0.295 1.380 0.465 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.520 2.205 0.960 2.635 ;
        RECT 1.520 2.205 2.380 2.635 ;
        RECT 2.600 2.035 2.925 2.465 ;
        RECT 0.085 1.865 2.085 2.035 ;
        RECT 0.085 1.495 0.395 1.865 ;
        RECT 0.085 0.825 0.255 1.495 ;
        RECT 1.405 0.825 1.575 1.325 ;
        RECT 1.915 0.995 2.085 1.865 ;
        RECT 2.255 1.455 2.925 2.035 ;
        RECT 3.450 1.875 3.830 2.635 ;
        RECT 2.255 0.825 2.470 1.455 ;
        RECT 0.085 0.430 0.345 0.825 ;
        RECT 0.645 0.085 0.825 0.825 ;
        RECT 1.405 0.655 2.470 0.825 ;
        RECT 1.560 0.085 1.925 0.465 ;
        RECT 2.140 0.255 2.470 0.655 ;
        RECT 2.695 0.735 3.890 0.905 ;
        RECT 2.695 0.365 2.945 0.735 ;
        RECT 3.165 0.085 3.335 0.555 ;
        RECT 3.555 0.270 3.890 0.735 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o21ba_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__o21ba_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o21ba_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 5.540 1.075 6.355 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 4.180 1.075 5.320 1.275 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.285 0.935 1.705 ;
        RECT 0.425 1.075 0.935 1.285 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.080 0.105 6.395 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.028500 ;
    PORT
      LAYER li1 ;
        RECT 1.155 1.445 2.425 1.705 ;
        RECT 1.155 0.910 1.705 1.445 ;
        RECT 1.155 0.725 2.375 0.910 ;
        RECT 1.155 0.255 1.485 0.725 ;
        RECT 2.045 0.255 2.375 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.085 2.045 0.435 2.465 ;
        RECT 0.635 2.215 1.015 2.635 ;
        RECT 1.575 2.215 1.955 2.635 ;
        RECT 2.515 2.215 2.895 2.635 ;
        RECT 0.085 1.875 2.815 2.045 ;
        RECT 0.085 1.455 0.435 1.875 ;
        RECT 2.645 1.615 2.815 1.875 ;
        RECT 3.115 1.965 3.285 2.465 ;
        RECT 3.550 2.135 3.800 2.635 ;
        RECT 4.035 2.295 5.265 2.465 ;
        RECT 4.035 2.135 4.325 2.295 ;
        RECT 4.585 1.965 4.830 2.125 ;
        RECT 3.115 1.795 4.830 1.965 ;
        RECT 0.085 0.855 0.255 1.455 ;
        RECT 2.645 1.445 3.205 1.615 ;
        RECT 1.875 1.080 2.815 1.250 ;
        RECT 0.085 0.265 0.545 0.855 ;
        RECT 0.765 0.085 0.935 0.905 ;
        RECT 2.645 0.895 2.815 1.080 ;
        RECT 2.985 1.245 3.205 1.445 ;
        RECT 2.985 1.075 3.435 1.245 ;
        RECT 3.745 0.895 3.935 1.795 ;
        RECT 4.585 1.445 4.830 1.795 ;
        RECT 5.095 1.665 5.265 2.295 ;
        RECT 5.435 1.835 5.815 2.635 ;
        RECT 6.035 1.665 6.310 2.465 ;
        RECT 5.095 1.455 6.310 1.665 ;
        RECT 2.645 0.645 3.935 0.895 ;
        RECT 4.155 0.725 6.310 0.905 ;
        RECT 1.705 0.085 1.875 0.555 ;
        RECT 4.155 0.475 4.405 0.725 ;
        RECT 2.565 0.085 2.895 0.475 ;
        RECT 3.105 0.255 4.405 0.475 ;
        RECT 4.625 0.085 4.795 0.555 ;
        RECT 4.965 0.255 5.345 0.725 ;
        RECT 5.565 0.085 5.735 0.555 ;
        RECT 5.905 0.265 6.310 0.725 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o21ba_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__o21bai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o21bai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.365 1.075 2.925 1.285 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.675 1.075 2.195 1.275 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.345 0.355 2.445 ;
        RECT 0.085 0.995 0.535 1.345 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.335 3.005 1.015 ;
        RECT 0.145 0.105 3.005 0.335 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.521500 ;
    PORT
      LAYER li1 ;
        RECT 1.635 1.625 2.155 2.465 ;
        RECT 1.235 1.445 2.155 1.625 ;
        RECT 1.235 0.255 1.455 1.445 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.525 1.705 0.850 2.210 ;
        RECT 1.070 1.875 1.400 2.635 ;
        RECT 0.525 1.535 1.065 1.705 ;
        RECT 2.470 1.535 3.060 2.635 ;
        RECT 0.770 0.995 1.065 1.535 ;
        RECT 0.770 0.825 0.940 0.995 ;
        RECT 0.085 0.085 0.360 0.825 ;
        RECT 0.675 0.495 0.940 0.825 ;
        RECT 1.640 0.735 2.915 0.905 ;
        RECT 1.640 0.255 1.970 0.735 ;
        RECT 2.195 0.085 2.365 0.555 ;
        RECT 2.535 0.270 2.915 0.735 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o21bai_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__o21bai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o21bai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 3.610 1.075 4.455 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.175 1.075 3.390 1.275 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.480 1.325 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.335 4.465 1.015 ;
        RECT 0.145 0.105 4.465 0.335 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.788000 ;
    PORT
      LAYER li1 ;
        RECT 1.185 1.615 1.355 2.465 ;
        RECT 2.655 1.615 2.900 2.125 ;
        RECT 1.185 1.445 2.900 1.615 ;
        RECT 1.510 0.645 2.005 1.445 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.180 1.665 0.350 1.915 ;
        RECT 0.635 1.875 0.965 2.635 ;
        RECT 1.620 1.795 1.870 2.635 ;
        RECT 2.105 2.295 3.335 2.465 ;
        RECT 2.105 1.795 2.435 2.295 ;
        RECT 3.165 1.665 3.335 2.295 ;
        RECT 3.505 1.835 3.885 2.635 ;
        RECT 4.105 1.665 4.380 2.465 ;
        RECT 0.180 1.495 0.915 1.665 ;
        RECT 0.650 1.245 0.915 1.495 ;
        RECT 3.165 1.455 4.380 1.665 ;
        RECT 0.650 1.075 1.340 1.245 ;
        RECT 0.180 0.085 0.350 0.825 ;
        RECT 0.650 0.445 0.820 1.075 ;
        RECT 1.060 0.475 1.340 0.905 ;
        RECT 2.225 0.725 4.380 0.905 ;
        RECT 2.225 0.475 2.475 0.725 ;
        RECT 1.060 0.255 2.475 0.475 ;
        RECT 2.695 0.085 2.865 0.555 ;
        RECT 3.035 0.255 3.415 0.725 ;
        RECT 3.635 0.085 3.805 0.555 ;
        RECT 3.975 0.265 4.380 0.725 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o21bai_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__o21bai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o21bai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 5.145 1.075 7.250 1.285 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 3.365 1.075 4.975 1.275 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.510 1.285 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.035 0.105 7.245 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.576000 ;
    PORT
      LAYER li1 ;
        RECT 1.035 1.625 1.375 2.465 ;
        RECT 2.065 1.625 2.315 2.465 ;
        RECT 3.575 1.625 3.825 2.125 ;
        RECT 4.515 1.625 4.765 2.125 ;
        RECT 1.035 1.455 4.765 1.625 ;
        RECT 2.695 1.445 4.765 1.455 ;
        RECT 2.695 1.075 3.195 1.445 ;
        RECT 2.695 0.815 2.925 1.075 ;
        RECT 1.520 0.645 2.925 0.815 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.360 2.805 ;
        RECT 0.145 1.625 0.475 2.435 ;
        RECT 0.695 1.795 0.865 2.635 ;
        RECT 1.595 1.795 1.845 2.635 ;
        RECT 2.535 1.795 2.785 2.635 ;
        RECT 3.025 2.295 5.235 2.465 ;
        RECT 3.025 1.795 3.355 2.295 ;
        RECT 4.045 1.795 4.295 2.295 ;
        RECT 4.985 1.625 5.235 2.295 ;
        RECT 5.455 1.795 5.705 2.635 ;
        RECT 5.925 1.625 6.175 2.465 ;
        RECT 6.395 1.795 6.645 2.635 ;
        RECT 6.865 1.625 7.115 2.465 ;
        RECT 0.145 1.455 0.850 1.625 ;
        RECT 4.985 1.455 7.115 1.625 ;
        RECT 0.680 1.285 0.850 1.455 ;
        RECT 0.680 1.075 2.525 1.285 ;
        RECT 0.680 0.895 0.945 1.075 ;
        RECT 0.225 0.085 0.395 0.895 ;
        RECT 0.565 0.290 0.945 0.895 ;
        RECT 3.145 0.725 7.155 0.905 ;
        RECT 3.145 0.475 3.395 0.725 ;
        RECT 1.180 0.305 3.395 0.475 ;
        RECT 3.615 0.085 3.785 0.555 ;
        RECT 3.955 0.255 4.335 0.725 ;
        RECT 4.555 0.085 4.725 0.555 ;
        RECT 4.895 0.255 5.275 0.725 ;
        RECT 5.495 0.085 5.665 0.555 ;
        RECT 5.835 0.255 6.215 0.725 ;
        RECT 6.435 0.085 6.605 0.555 ;
        RECT 6.775 0.255 7.155 0.725 ;
        RECT 0.000 -0.085 7.360 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o21bai_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__o22a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o22a_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.835 1.075 3.310 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.325 2.665 2.405 ;
        RECT 2.335 1.075 2.665 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.075 1.535 1.325 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.730 1.075 2.155 1.325 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.435 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.472000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.365 0.365 2.465 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.605 1.875 1.360 2.635 ;
        RECT 1.805 1.705 2.275 2.465 ;
        RECT 0.535 1.495 2.275 1.705 ;
        RECT 0.535 0.895 0.860 1.495 ;
        RECT 2.985 1.455 3.540 2.635 ;
        RECT 0.535 0.715 1.805 0.895 ;
        RECT 1.440 0.645 1.805 0.715 ;
        RECT 2.065 0.695 3.355 0.865 ;
        RECT 0.615 0.085 0.785 0.545 ;
        RECT 2.065 0.475 2.395 0.695 ;
        RECT 1.055 0.295 2.395 0.475 ;
        RECT 2.625 0.085 2.795 0.525 ;
        RECT 2.965 0.280 3.355 0.695 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o22a_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__o22a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o22a_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 3.345 1.075 3.705 1.615 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.905 1.275 3.175 2.405 ;
        RECT 2.795 1.075 3.175 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.525 1.075 1.890 1.275 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.110 1.075 2.625 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.015 0.105 3.975 1.015 ;
        RECT 0.130 -0.085 0.300 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.491500 ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.365 0.855 2.465 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.115 1.445 0.365 2.635 ;
        RECT 1.095 1.875 1.895 2.635 ;
        RECT 2.340 1.705 2.695 2.465 ;
        RECT 3.570 1.795 3.890 2.635 ;
        RECT 1.075 1.455 2.695 1.705 ;
        RECT 1.075 0.895 1.355 1.455 ;
        RECT 0.185 0.085 0.355 0.885 ;
        RECT 1.075 0.715 2.365 0.895 ;
        RECT 1.950 0.645 2.365 0.715 ;
        RECT 2.590 0.695 3.890 0.865 ;
        RECT 1.125 0.085 1.305 0.545 ;
        RECT 2.590 0.475 2.930 0.695 ;
        RECT 1.565 0.295 2.930 0.475 ;
        RECT 3.195 0.085 3.365 0.525 ;
        RECT 3.555 0.280 3.890 0.695 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o22a_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__o22a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o22a_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.900 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 4.710 1.445 6.285 1.615 ;
        RECT 4.710 1.075 5.130 1.445 ;
        RECT 6.075 1.275 6.285 1.445 ;
        RECT 6.075 1.075 6.815 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 5.350 1.075 5.905 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.620 1.445 4.540 1.615 ;
        RECT 2.620 1.075 3.180 1.445 ;
        RECT 4.200 1.075 4.540 1.445 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 3.350 1.075 4.030 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.900 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.070 0.105 6.840 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.090 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.900 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.028500 ;
    PORT
      LAYER li1 ;
        RECT 0.690 1.615 0.940 2.465 ;
        RECT 1.630 1.615 1.880 2.465 ;
        RECT 0.085 1.445 1.880 1.615 ;
        RECT 0.085 0.905 0.370 1.445 ;
        RECT 0.085 0.725 1.920 0.905 ;
        RECT 0.600 0.265 0.980 0.725 ;
        RECT 1.540 0.255 1.920 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.900 2.805 ;
        RECT 0.220 1.825 0.470 2.635 ;
        RECT 1.160 1.795 1.410 2.635 ;
        RECT 2.100 2.125 2.870 2.635 ;
        RECT 3.090 2.295 4.280 2.465 ;
        RECT 3.090 2.125 3.340 2.295 ;
        RECT 4.030 2.125 4.280 2.295 ;
        RECT 4.500 2.125 4.830 2.635 ;
        RECT 5.050 2.295 6.240 2.465 ;
        RECT 5.050 2.125 5.300 2.295 ;
        RECT 3.560 1.955 3.810 2.125 ;
        RECT 5.520 1.955 5.770 2.125 ;
        RECT 2.100 1.785 5.770 1.955 ;
        RECT 5.990 1.785 6.240 2.295 ;
        RECT 2.100 1.275 2.430 1.785 ;
        RECT 6.505 1.455 6.710 2.635 ;
        RECT 0.540 1.075 2.430 1.275 ;
        RECT 2.140 0.905 2.430 1.075 ;
        RECT 2.140 0.735 4.320 0.905 ;
        RECT 2.615 0.645 4.320 0.735 ;
        RECT 4.540 0.735 6.750 0.905 ;
        RECT 0.260 0.085 0.430 0.555 ;
        RECT 1.200 0.085 1.370 0.555 ;
        RECT 2.140 0.085 2.310 0.555 ;
        RECT 4.540 0.475 4.870 0.735 ;
        RECT 5.430 0.725 6.750 0.735 ;
        RECT 2.580 0.255 4.870 0.475 ;
        RECT 5.090 0.085 5.260 0.555 ;
        RECT 5.430 0.255 5.810 0.725 ;
        RECT 6.030 0.085 6.200 0.555 ;
        RECT 6.370 0.255 6.750 0.725 ;
        RECT 0.000 -0.085 6.900 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o22a_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__o22ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o22ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.150 1.075 2.660 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.920 1.615 2.170 2.405 ;
        RECT 1.750 1.445 2.170 1.615 ;
        RECT 1.750 1.245 1.980 1.445 ;
        RECT 1.565 1.075 1.980 1.245 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.665 0.325 1.990 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.050 0.995 1.350 1.665 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.740 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.816750 ;
    PORT
      LAYER li1 ;
        RECT 1.130 2.045 1.680 2.465 ;
        RECT 0.495 1.835 1.680 2.045 ;
        RECT 0.495 0.825 0.790 1.835 ;
        RECT 0.495 0.645 0.895 0.825 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.135 2.175 0.345 2.635 ;
        RECT 2.340 1.455 2.660 2.635 ;
        RECT 1.460 0.825 2.660 0.865 ;
        RECT 1.290 0.695 2.660 0.825 ;
        RECT 1.290 0.475 1.620 0.695 ;
        RECT 0.085 0.295 1.620 0.475 ;
        RECT 1.890 0.085 2.060 0.525 ;
        RECT 2.270 0.280 2.660 0.695 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o22ai_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__o22ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o22ai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 3.765 1.075 4.565 1.285 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.835 1.075 3.555 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.200 1.075 1.115 1.285 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 1.325 1.075 2.125 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.855 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.061000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.625 1.815 2.125 ;
        RECT 3.065 1.625 3.315 2.125 ;
        RECT 1.565 1.445 3.315 1.625 ;
        RECT 2.405 0.905 2.645 1.445 ;
        RECT 0.535 0.645 2.645 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.060 2.805 ;
        RECT 0.150 1.625 0.405 2.465 ;
        RECT 0.625 1.795 0.875 2.635 ;
        RECT 1.095 2.295 2.285 2.465 ;
        RECT 1.095 1.625 1.345 2.295 ;
        RECT 2.035 1.795 2.285 2.295 ;
        RECT 2.595 2.295 3.785 2.465 ;
        RECT 2.595 1.795 2.845 2.295 ;
        RECT 0.150 1.455 1.345 1.625 ;
        RECT 3.535 1.625 3.785 2.295 ;
        RECT 4.005 1.795 4.255 2.635 ;
        RECT 4.475 1.625 4.730 2.465 ;
        RECT 3.535 1.455 4.730 1.625 ;
        RECT 0.090 0.475 0.365 0.905 ;
        RECT 2.815 0.725 4.765 0.905 ;
        RECT 2.815 0.475 2.985 0.725 ;
        RECT 0.090 0.305 2.985 0.475 ;
        RECT 3.155 0.085 3.325 0.555 ;
        RECT 3.495 0.255 3.825 0.725 ;
        RECT 4.045 0.085 4.215 0.555 ;
        RECT 4.385 0.255 4.765 0.725 ;
        RECT 0.000 -0.085 5.060 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o22ai_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__o22ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o22ai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.280 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 1.250 1.445 4.030 1.615 ;
        RECT 1.250 1.275 1.565 1.445 ;
        RECT 0.085 1.075 1.565 1.275 ;
        RECT 3.625 1.075 4.030 1.445 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 1.835 1.075 3.445 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 4.745 1.445 7.735 1.615 ;
        RECT 4.745 0.995 5.490 1.445 ;
        RECT 7.465 0.995 7.735 1.445 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 5.660 1.075 7.160 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.280 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.035 0.105 8.115 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.470 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.280 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.959500 ;
    PORT
      LAYER li1 ;
        RECT 1.955 1.955 2.295 2.125 ;
        RECT 2.985 1.955 3.235 2.125 ;
        RECT 5.855 1.955 6.105 2.125 ;
        RECT 6.795 1.955 7.045 2.125 ;
        RECT 1.955 1.785 4.370 1.955 ;
        RECT 5.855 1.785 8.170 1.955 ;
        RECT 4.200 1.615 4.370 1.785 ;
        RECT 4.200 1.445 4.575 1.615 ;
        RECT 4.355 0.820 4.575 1.445 ;
        RECT 7.905 0.820 8.170 1.785 ;
        RECT 4.355 0.645 8.170 0.820 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.280 2.805 ;
        RECT 0.165 1.445 0.415 2.635 ;
        RECT 0.635 1.955 0.885 2.465 ;
        RECT 1.105 2.125 1.355 2.635 ;
        RECT 1.575 2.295 3.745 2.465 ;
        RECT 1.575 1.955 1.785 2.295 ;
        RECT 2.515 2.125 2.765 2.295 ;
        RECT 3.455 2.125 3.745 2.295 ;
        RECT 3.965 2.125 4.185 2.635 ;
        RECT 4.355 2.125 4.710 2.465 ;
        RECT 4.925 2.125 5.165 2.635 ;
        RECT 5.385 2.295 7.515 2.465 ;
        RECT 0.635 1.785 1.785 1.955 ;
        RECT 4.540 1.955 4.710 2.125 ;
        RECT 5.385 1.955 5.635 2.295 ;
        RECT 6.325 2.125 6.575 2.295 ;
        RECT 7.265 2.135 7.515 2.295 ;
        RECT 7.735 2.125 8.015 2.635 ;
        RECT 4.540 1.785 5.635 1.955 ;
        RECT 0.635 1.445 0.885 1.785 ;
        RECT 0.125 0.735 4.185 0.905 ;
        RECT 0.125 0.725 1.395 0.735 ;
        RECT 0.125 0.255 0.455 0.725 ;
        RECT 0.675 0.085 0.845 0.555 ;
        RECT 1.015 0.255 1.395 0.725 ;
        RECT 1.955 0.725 3.275 0.735 ;
        RECT 1.615 0.085 1.785 0.555 ;
        RECT 1.955 0.255 2.335 0.725 ;
        RECT 2.555 0.085 2.725 0.555 ;
        RECT 2.895 0.255 3.275 0.725 ;
        RECT 3.495 0.085 3.665 0.555 ;
        RECT 3.835 0.475 4.185 0.735 ;
        RECT 3.835 0.255 8.045 0.475 ;
        RECT 0.000 -0.085 8.280 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o22ai_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__o31ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o31ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 0.435 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.075 1.105 2.465 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.455 1.325 1.695 2.405 ;
        RECT 1.315 1.075 1.695 1.325 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.325 0.995 2.650 1.325 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.655 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.833500 ;
    PORT
      LAYER li1 ;
        RECT 1.885 0.825 2.155 2.465 ;
        RECT 1.885 0.260 2.495 0.825 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT -0.015 2.635 2.760 2.805 ;
        RECT 0.085 1.495 0.420 2.635 ;
        RECT 2.355 1.495 2.525 2.635 ;
        RECT 0.175 0.085 0.345 0.905 ;
        RECT 0.515 0.735 1.715 0.905 ;
        RECT 0.515 0.255 0.895 0.735 ;
        RECT 1.125 0.085 1.295 0.565 ;
        RECT 1.465 0.460 1.715 0.735 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o31ai_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__o31ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o31ai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.055 1.310 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 1.500 1.055 2.420 1.325 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.700 1.055 3.555 1.325 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 4.630 0.755 4.970 1.325 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.010 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.136000 ;
    PORT
      LAYER li1 ;
        RECT 2.585 1.665 2.915 2.125 ;
        RECT 3.475 1.665 3.855 2.465 ;
        RECT 4.625 1.665 4.965 2.465 ;
        RECT 2.585 1.495 4.965 1.665 ;
        RECT 4.075 0.595 4.455 1.495 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.060 2.805 ;
        RECT 0.090 1.665 0.445 2.465 ;
        RECT 0.665 1.835 0.835 2.635 ;
        RECT 1.005 1.665 1.385 2.465 ;
        RECT 1.605 2.295 3.305 2.465 ;
        RECT 1.605 1.835 1.775 2.295 ;
        RECT 1.945 1.665 2.325 2.125 ;
        RECT 3.135 1.835 3.305 2.295 ;
        RECT 4.075 1.835 4.405 2.635 ;
        RECT 0.090 1.495 2.325 1.665 ;
        RECT 0.090 0.715 3.855 0.885 ;
        RECT 0.090 0.255 0.445 0.715 ;
        RECT 0.665 0.085 0.835 0.545 ;
        RECT 1.005 0.255 1.385 0.715 ;
        RECT 1.605 0.085 2.165 0.545 ;
        RECT 2.425 0.255 2.755 0.715 ;
        RECT 2.925 0.085 3.305 0.545 ;
        RECT 3.475 0.425 3.855 0.715 ;
        RECT 4.630 0.425 4.965 0.585 ;
        RECT 3.475 0.255 4.965 0.425 ;
        RECT 0.000 -0.085 5.060 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o31ai_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__o31ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o31ai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.740 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.055 1.930 1.425 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 2.150 1.055 4.005 1.425 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 4.175 1.055 6.590 1.275 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 7.165 1.055 8.585 1.275 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.740 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.025 0.105 8.640 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.930 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.740 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.851000 ;
    PORT
      LAYER li1 ;
        RECT 6.420 1.695 6.590 2.465 ;
        RECT 7.360 1.695 7.530 2.465 ;
        RECT 8.300 1.695 8.625 2.465 ;
        RECT 4.175 1.445 8.625 1.695 ;
        RECT 6.760 0.885 6.995 1.445 ;
        RECT 6.760 0.645 8.080 0.885 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.740 2.805 ;
        RECT 0.090 1.895 0.445 2.465 ;
        RECT 0.665 2.065 0.835 2.635 ;
        RECT 1.005 1.895 1.385 2.465 ;
        RECT 1.605 2.065 1.775 2.635 ;
        RECT 1.945 2.205 4.285 2.465 ;
        RECT 1.945 1.895 2.325 2.205 ;
        RECT 0.090 1.595 2.325 1.895 ;
        RECT 2.545 1.765 2.715 2.035 ;
        RECT 2.885 1.935 3.265 2.205 ;
        RECT 4.530 2.035 6.200 2.465 ;
        RECT 3.485 1.865 6.200 2.035 ;
        RECT 6.760 1.890 7.140 2.635 ;
        RECT 7.700 1.890 8.080 2.635 ;
        RECT 3.485 1.765 4.005 1.865 ;
        RECT 2.545 1.595 4.005 1.765 ;
        RECT 0.090 0.715 6.590 0.885 ;
        RECT 0.090 0.255 0.445 0.715 ;
        RECT 0.665 0.085 0.835 0.545 ;
        RECT 1.005 0.255 1.385 0.715 ;
        RECT 1.605 0.085 1.775 0.545 ;
        RECT 1.945 0.255 2.325 0.715 ;
        RECT 2.545 0.085 2.715 0.545 ;
        RECT 2.885 0.255 3.265 0.715 ;
        RECT 3.485 0.085 3.655 0.545 ;
        RECT 3.825 0.255 4.205 0.715 ;
        RECT 4.445 0.085 5.140 0.545 ;
        RECT 5.360 0.395 5.530 0.715 ;
        RECT 5.790 0.085 6.160 0.545 ;
        RECT 6.420 0.475 6.590 0.715 ;
        RECT 8.300 0.475 8.585 0.885 ;
        RECT 6.420 0.255 8.585 0.475 ;
        RECT 0.000 -0.085 8.740 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o31ai_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__o32ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o32ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.395 0.995 2.990 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.915 0.995 2.205 2.465 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.475 0.995 1.745 1.615 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.685 0.360 1.325 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.920 0.995 1.305 1.615 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.185 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.758750 ;
    PORT
      LAYER li1 ;
        RECT 0.530 1.785 1.530 2.465 ;
        RECT 0.530 0.825 0.750 1.785 ;
        RECT 0.530 0.655 0.895 0.825 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.090 1.495 0.360 2.635 ;
        RECT 2.785 1.495 3.135 2.635 ;
        RECT 1.065 0.655 2.555 0.825 ;
        RECT 1.065 0.485 1.440 0.655 ;
        RECT 0.085 0.255 1.440 0.485 ;
        RECT 1.645 0.085 1.975 0.485 ;
        RECT 2.385 0.375 2.555 0.655 ;
        RECT 2.725 0.085 3.095 0.825 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o32ai_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__o32ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o32ai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 5.200 1.075 6.295 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 3.720 1.075 4.930 1.325 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.655 1.075 3.365 1.325 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.075 1.815 1.325 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 0.895 1.325 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 6.395 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.061000 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.665 0.895 2.095 ;
        RECT 3.025 1.665 3.405 2.085 ;
        RECT 0.515 1.495 3.405 1.665 ;
        RECT 1.985 1.105 2.370 1.495 ;
        RECT 1.985 0.905 2.245 1.105 ;
        RECT 0.515 0.655 2.245 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.090 2.295 1.365 2.465 ;
        RECT 0.090 1.495 0.345 2.295 ;
        RECT 1.115 2.005 1.365 2.295 ;
        RECT 1.585 2.175 1.755 2.635 ;
        RECT 1.925 2.005 2.305 2.455 ;
        RECT 1.115 1.835 2.305 2.005 ;
        RECT 2.585 2.255 4.835 2.445 ;
        RECT 2.585 1.835 2.835 2.255 ;
        RECT 3.625 1.495 3.795 2.255 ;
        RECT 4.015 1.665 4.345 2.085 ;
        RECT 4.585 1.835 4.835 2.255 ;
        RECT 5.070 1.835 5.275 2.635 ;
        RECT 5.495 1.665 5.825 2.460 ;
        RECT 4.015 1.495 5.825 1.665 ;
        RECT 6.045 1.495 6.265 2.635 ;
        RECT 0.090 0.485 0.345 0.905 ;
        RECT 2.485 0.715 6.305 0.905 ;
        RECT 2.485 0.485 2.655 0.715 ;
        RECT 0.090 0.255 2.655 0.485 ;
        RECT 2.870 0.085 3.250 0.545 ;
        RECT 3.435 0.255 3.815 0.715 ;
        RECT 4.035 0.085 4.205 0.545 ;
        RECT 4.505 0.255 5.175 0.715 ;
        RECT 5.355 0.085 5.735 0.545 ;
        RECT 5.975 0.255 6.305 0.715 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o32ai_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__o32ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o32ai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.040 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 9.090 1.075 10.925 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 6.520 1.075 8.010 1.275 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 4.170 1.075 5.980 1.275 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 2.405 1.075 3.940 1.275 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.110 1.075 1.835 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.040 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 11.015 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 11.230 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.040 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.024500 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.665 0.895 2.085 ;
        RECT 1.455 1.665 1.850 2.085 ;
        RECT 4.860 1.665 5.190 2.085 ;
        RECT 5.750 1.665 6.130 2.085 ;
        RECT 0.515 1.495 6.130 1.665 ;
        RECT 2.055 0.905 2.235 1.495 ;
        RECT 0.515 0.655 3.730 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 11.040 2.805 ;
        RECT 0.090 2.255 2.240 2.465 ;
        RECT 0.090 1.495 0.345 2.255 ;
        RECT 1.115 1.835 1.285 2.255 ;
        RECT 2.070 2.005 2.240 2.255 ;
        RECT 2.410 2.175 2.790 2.635 ;
        RECT 3.010 2.005 3.180 2.425 ;
        RECT 3.350 2.175 3.730 2.635 ;
        RECT 3.950 2.005 4.200 2.465 ;
        RECT 2.070 1.835 4.200 2.005 ;
        RECT 4.390 2.255 8.480 2.465 ;
        RECT 4.390 1.835 4.640 2.255 ;
        RECT 5.410 1.835 5.580 2.255 ;
        RECT 6.350 1.835 6.520 2.255 ;
        RECT 6.690 1.665 7.070 2.085 ;
        RECT 7.290 1.835 7.460 2.255 ;
        RECT 7.630 1.665 8.010 2.085 ;
        RECT 8.230 1.835 8.480 2.255 ;
        RECT 8.670 1.835 8.920 2.635 ;
        RECT 9.090 1.665 9.470 2.465 ;
        RECT 9.690 1.835 9.860 2.635 ;
        RECT 10.030 1.665 10.410 2.465 ;
        RECT 6.690 1.495 10.410 1.665 ;
        RECT 10.675 1.495 10.925 2.635 ;
        RECT 0.090 0.465 0.345 0.905 ;
        RECT 3.950 0.735 10.925 0.905 ;
        RECT 3.950 0.465 4.200 0.735 ;
        RECT 0.090 0.255 4.200 0.465 ;
        RECT 4.420 0.085 4.590 0.545 ;
        RECT 4.760 0.255 5.140 0.735 ;
        RECT 5.360 0.085 5.690 0.545 ;
        RECT 5.910 0.255 6.580 0.735 ;
        RECT 6.820 0.085 6.990 0.545 ;
        RECT 7.160 0.255 7.540 0.735 ;
        RECT 7.760 0.085 7.930 0.545 ;
        RECT 8.100 0.255 8.840 0.735 ;
        RECT 9.220 0.085 9.390 0.545 ;
        RECT 9.560 0.255 9.940 0.735 ;
        RECT 10.160 0.085 10.375 0.545 ;
        RECT 10.545 0.255 10.925 0.735 ;
        RECT 0.000 -0.085 11.040 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o32ai_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__o211a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o211a_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.350 1.075 1.815 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.985 1.075 2.370 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.540 1.075 3.080 1.275 ;
        RECT 2.815 0.435 3.080 1.075 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 3.640 1.075 4.005 1.325 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.890 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.495 0.425 2.465 ;
        RECT 0.085 0.885 0.260 1.495 ;
        RECT 0.085 0.255 0.425 0.885 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.645 1.495 0.815 2.635 ;
        RECT 1.085 1.835 1.335 2.635 ;
        RECT 2.085 1.665 2.465 2.465 ;
        RECT 2.760 1.835 3.090 2.635 ;
        RECT 3.470 1.665 3.800 2.465 ;
        RECT 1.005 1.495 3.800 1.665 ;
        RECT 1.005 1.245 1.175 1.495 ;
        RECT 0.430 1.075 1.175 1.245 ;
        RECT 0.645 0.085 0.895 0.885 ;
        RECT 1.085 0.735 2.410 0.905 ;
        RECT 1.085 0.255 1.415 0.735 ;
        RECT 1.635 0.085 1.860 0.545 ;
        RECT 2.030 0.255 2.410 0.735 ;
        RECT 3.250 0.865 3.470 1.495 ;
        RECT 3.250 0.255 3.800 0.865 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o211a_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__o211a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o211a_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.165 0.995 2.675 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.505 0.995 1.945 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.930 0.995 1.310 1.325 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.360 1.325 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.120 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.534000 ;
    PORT
      LAYER li1 ;
        RECT 3.085 2.075 3.275 2.465 ;
        RECT 3.085 1.905 4.035 2.075 ;
        RECT 3.765 0.785 4.035 1.905 ;
        RECT 2.945 0.615 4.035 0.785 ;
        RECT 2.945 0.255 3.325 0.615 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.090 1.765 0.355 2.465 ;
        RECT 0.525 1.935 0.905 2.635 ;
        RECT 1.125 1.765 1.820 2.465 ;
        RECT 2.375 1.935 2.855 2.635 ;
        RECT 3.445 2.255 3.825 2.635 ;
        RECT 0.090 1.735 1.820 1.765 ;
        RECT 0.090 1.510 3.025 1.735 ;
        RECT 0.530 0.825 0.760 1.510 ;
        RECT 2.855 1.325 3.025 1.510 ;
        RECT 2.855 0.995 3.565 1.325 ;
        RECT 0.095 0.425 0.760 0.825 ;
        RECT 0.930 0.635 2.375 0.825 ;
        RECT 0.095 0.255 0.430 0.425 ;
        RECT 1.535 0.085 1.870 0.465 ;
        RECT 2.540 0.085 2.775 0.525 ;
        RECT 3.545 0.085 3.875 0.445 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o211a_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__o211a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o211a_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.900 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 4.825 1.495 6.815 1.685 ;
        RECT 4.825 1.035 5.155 1.495 ;
        RECT 6.300 1.035 6.815 1.495 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 5.340 1.035 6.115 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.790 1.445 4.600 1.685 ;
        RECT 2.790 0.995 3.085 1.445 ;
        RECT 4.270 1.035 4.600 1.445 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 3.255 1.035 4.090 1.275 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.900 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 6.895 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.090 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.900 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.016000 ;
    PORT
      LAYER li1 ;
        RECT 1.080 1.700 1.260 2.465 ;
        RECT 2.040 1.700 2.230 2.465 ;
        RECT 0.085 1.435 2.230 1.700 ;
        RECT 0.085 0.805 0.365 1.435 ;
        RECT 0.085 0.635 1.755 0.805 ;
        RECT 0.645 0.615 1.755 0.635 ;
        RECT 0.645 0.255 0.815 0.615 ;
        RECT 1.585 0.255 1.755 0.615 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.900 2.805 ;
        RECT 0.480 1.870 0.860 2.635 ;
        RECT 1.440 1.870 1.820 2.635 ;
        RECT 2.400 2.200 2.780 2.635 ;
        RECT 3.000 2.025 3.360 2.465 ;
        RECT 3.535 2.195 3.915 2.635 ;
        RECT 4.085 2.025 4.415 2.465 ;
        RECT 4.595 2.195 4.860 2.635 ;
        RECT 5.465 2.025 5.845 2.465 ;
        RECT 2.400 1.855 5.845 2.025 ;
        RECT 6.425 1.915 6.805 2.635 ;
        RECT 2.400 1.265 2.620 1.855 ;
        RECT 0.535 1.065 2.620 1.265 ;
        RECT 2.400 0.815 2.620 1.065 ;
        RECT 2.400 0.635 3.820 0.815 ;
        RECT 4.475 0.695 6.805 0.865 ;
        RECT 4.475 0.465 4.805 0.695 ;
        RECT 0.095 0.085 0.425 0.465 ;
        RECT 1.035 0.085 1.365 0.445 ;
        RECT 1.925 0.085 2.340 0.465 ;
        RECT 2.580 0.255 4.805 0.465 ;
        RECT 4.980 0.085 5.295 0.525 ;
        RECT 5.465 0.255 5.845 0.695 ;
        RECT 6.065 0.085 6.255 0.525 ;
        RECT 6.425 0.255 6.805 0.695 ;
        RECT 0.000 -0.085 6.900 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o211a_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__o211ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o211ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.395 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.565 1.325 0.825 2.250 ;
        RECT 0.565 0.995 1.080 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.495 1.345 1.745 1.615 ;
        RECT 1.420 0.995 1.745 1.345 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.915 1.020 2.270 1.615 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.755 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.297000 ;
    PORT
      LAYER li1 ;
        RECT 0.995 2.045 1.325 2.445 ;
        RECT 2.075 2.045 2.675 2.465 ;
        RECT 0.995 1.815 2.675 2.045 ;
        RECT 0.995 1.595 1.325 1.815 ;
        RECT 2.440 0.825 2.675 1.815 ;
        RECT 1.725 0.255 2.675 0.825 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.095 1.495 0.395 2.635 ;
        RECT 1.540 2.275 1.870 2.635 ;
        RECT 0.095 0.615 1.450 0.825 ;
        RECT 0.095 0.255 0.400 0.615 ;
        RECT 0.570 0.085 0.900 0.445 ;
        RECT 1.070 0.255 1.450 0.615 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o211ai_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__o211ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o211ai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 3.805 1.075 4.915 1.295 ;
        RECT 4.465 0.765 4.915 1.075 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.670 1.075 3.635 1.355 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 1.215 1.075 2.210 1.365 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.375 1.970 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.980 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.114500 ;
    PORT
      LAYER li1 ;
        RECT 0.545 1.710 0.855 2.465 ;
        RECT 1.625 1.710 1.815 2.465 ;
        RECT 3.025 1.710 3.405 2.125 ;
        RECT 0.545 1.540 3.405 1.710 ;
        RECT 0.545 0.670 0.925 1.540 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.060 2.805 ;
        RECT 0.115 2.175 0.375 2.635 ;
        RECT 1.025 1.915 1.405 2.635 ;
        RECT 1.985 1.915 2.365 2.635 ;
        RECT 2.595 2.295 3.815 2.465 ;
        RECT 2.595 2.100 2.855 2.295 ;
        RECT 3.625 1.695 3.815 2.295 ;
        RECT 3.985 1.865 4.365 2.635 ;
        RECT 4.585 1.695 4.845 2.465 ;
        RECT 3.625 1.525 4.845 1.695 ;
        RECT 1.145 0.465 1.335 0.890 ;
        RECT 1.505 0.635 4.295 0.845 ;
        RECT 4.105 0.515 4.295 0.635 ;
        RECT 1.145 0.445 2.365 0.465 ;
        RECT 0.095 0.255 2.365 0.445 ;
        RECT 2.595 0.085 2.925 0.445 ;
        RECT 3.525 0.085 3.905 0.445 ;
        RECT 4.465 0.085 4.870 0.445 ;
        RECT 0.000 -0.085 5.060 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o211ai_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__o211ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o211ai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.740 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 1.015 1.515 4.030 1.685 ;
        RECT 1.015 1.330 1.560 1.515 ;
        RECT 0.400 1.075 1.560 1.330 ;
        RECT 3.700 0.995 4.030 1.515 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 1.855 1.075 3.530 1.345 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 4.710 1.515 7.800 1.685 ;
        RECT 4.710 1.410 5.525 1.515 ;
        RECT 4.200 0.995 5.525 1.410 ;
        RECT 7.580 0.995 7.800 1.515 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 5.970 1.075 7.140 1.345 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.740 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 8.375 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.930 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.740 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.218500 ;
    PORT
      LAYER li1 ;
        RECT 1.955 2.025 3.820 2.105 ;
        RECT 4.495 2.025 8.480 2.105 ;
        RECT 1.955 1.855 8.480 2.025 ;
        RECT 7.980 1.340 8.480 1.855 ;
        RECT 7.980 0.825 8.160 1.340 ;
        RECT 7.265 0.655 8.160 0.825 ;
        RECT 7.265 0.450 7.485 0.655 ;
        RECT 5.830 0.270 7.485 0.450 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.740 2.805 ;
        RECT 0.090 1.665 0.385 2.635 ;
        RECT 1.005 2.275 1.385 2.635 ;
        RECT 1.605 2.275 3.785 2.465 ;
        RECT 0.605 2.105 0.825 2.190 ;
        RECT 1.605 2.105 1.785 2.275 ;
        RECT 4.015 2.195 4.285 2.635 ;
        RECT 4.885 2.275 5.265 2.635 ;
        RECT 5.830 2.275 6.210 2.635 ;
        RECT 6.770 2.275 7.155 2.635 ;
        RECT 8.155 2.275 8.485 2.635 ;
        RECT 0.605 1.935 1.785 2.105 ;
        RECT 0.605 1.860 0.825 1.935 ;
        RECT 0.155 0.795 3.480 0.905 ;
        RECT 0.155 0.625 4.235 0.795 ;
        RECT 4.405 0.635 6.870 0.815 ;
        RECT 0.155 0.535 0.355 0.625 ;
        RECT 0.525 0.085 0.905 0.445 ;
        RECT 1.125 0.425 1.340 0.625 ;
        RECT 4.005 0.455 4.235 0.625 ;
        RECT 8.320 0.480 8.490 0.595 ;
        RECT 1.535 0.085 1.865 0.455 ;
        RECT 2.445 0.085 2.825 0.445 ;
        RECT 3.405 0.085 3.785 0.445 ;
        RECT 4.005 0.255 5.470 0.455 ;
        RECT 7.730 0.310 8.490 0.480 ;
        RECT 0.000 -0.085 8.740 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 1.170 0.425 1.340 0.595 ;
        RECT 8.320 0.425 8.490 0.595 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
      LAYER met1 ;
        RECT 1.110 0.580 1.400 0.625 ;
        RECT 8.260 0.580 8.550 0.625 ;
        RECT 1.110 0.440 8.550 0.580 ;
        RECT 1.110 0.395 1.400 0.440 ;
        RECT 8.260 0.395 8.550 0.440 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o211ai_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__o221a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o221a_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.815 1.075 3.145 1.285 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.980 1.255 2.315 1.705 ;
        RECT 1.980 0.985 2.615 1.255 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.925 0.985 1.235 1.325 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.405 0.985 1.790 1.705 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.415 1.285 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.080 0.105 3.935 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.504500 ;
    PORT
      LAYER li1 ;
        RECT 3.465 1.875 4.030 2.465 ;
        RECT 3.715 0.825 4.030 1.875 ;
        RECT 3.445 0.265 4.030 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.085 1.720 0.365 2.465 ;
        RECT 0.560 2.085 0.860 2.635 ;
        RECT 1.500 2.045 2.355 2.465 ;
        RECT 1.030 1.875 2.745 2.045 ;
        RECT 1.030 1.720 1.235 1.875 ;
        RECT 0.085 1.495 1.235 1.720 ;
        RECT 2.575 1.625 2.745 1.875 ;
        RECT 2.915 1.795 3.295 2.635 ;
        RECT 0.085 1.455 0.755 1.495 ;
        RECT 2.575 1.455 3.545 1.625 ;
        RECT 0.585 0.825 0.755 1.455 ;
        RECT 3.375 0.995 3.545 1.455 ;
        RECT 0.170 0.645 0.755 0.825 ;
        RECT 1.035 0.645 2.935 0.815 ;
        RECT 0.170 0.255 0.500 0.645 ;
        RECT 0.700 0.305 1.905 0.475 ;
        RECT 2.085 0.085 2.425 0.475 ;
        RECT 2.605 0.270 2.935 0.645 ;
        RECT 3.105 0.085 3.275 0.640 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o221a_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__o221a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o221a_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.835 1.075 3.325 1.285 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.235 1.075 2.615 1.705 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.935 1.075 1.330 1.275 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.520 1.075 1.905 1.705 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.345 1.325 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.060 0.105 4.485 1.015 ;
        RECT 0.120 -0.085 0.290 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.530500 ;
    PORT
      LAYER li1 ;
        RECT 3.545 2.045 3.845 2.465 ;
        RECT 3.545 1.875 4.490 2.045 ;
        RECT 4.180 0.905 4.490 1.875 ;
        RECT 3.545 0.735 4.490 0.905 ;
        RECT 3.545 0.265 3.925 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.250 1.670 0.580 2.465 ;
        RECT 0.800 1.850 1.010 2.635 ;
        RECT 1.700 2.045 2.455 2.465 ;
        RECT 1.180 1.875 2.965 2.045 ;
        RECT 1.180 1.670 1.350 1.875 ;
        RECT 0.250 1.495 1.350 1.670 ;
        RECT 0.545 1.445 1.350 1.495 ;
        RECT 2.795 1.625 2.965 1.875 ;
        RECT 3.145 1.795 3.375 2.635 ;
        RECT 4.015 2.215 4.405 2.635 ;
        RECT 2.795 1.455 3.715 1.625 ;
        RECT 0.545 0.805 0.765 1.445 ;
        RECT 3.495 1.285 3.715 1.455 ;
        RECT 3.495 1.075 3.875 1.285 ;
        RECT 0.170 0.635 0.765 0.805 ;
        RECT 1.135 0.735 2.985 0.905 ;
        RECT 1.135 0.645 1.570 0.735 ;
        RECT 0.170 0.255 0.500 0.635 ;
        RECT 0.670 0.295 2.005 0.465 ;
        RECT 2.265 0.085 2.435 0.555 ;
        RECT 2.605 0.270 2.985 0.735 ;
        RECT 3.205 0.085 3.375 0.905 ;
        RECT 4.145 0.085 4.315 0.565 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o221a_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__o221a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o221a_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.820 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 3.305 1.445 5.225 1.615 ;
        RECT 3.305 1.075 3.955 1.445 ;
        RECT 4.975 1.275 5.225 1.445 ;
        RECT 4.975 1.075 5.535 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 4.125 1.075 4.755 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.445 3.045 1.615 ;
        RECT 1.065 1.075 1.730 1.445 ;
        RECT 2.665 1.075 3.045 1.445 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 1.950 1.075 2.495 1.275 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 0.440 1.275 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.820 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 7.615 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.010 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.820 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.028500 ;
    PORT
      LAYER li1 ;
        RECT 5.865 1.955 6.075 2.465 ;
        RECT 5.865 1.785 6.500 1.955 ;
        RECT 6.330 1.615 6.500 1.785 ;
        RECT 6.765 1.615 7.015 2.465 ;
        RECT 6.330 1.445 7.710 1.615 ;
        RECT 7.365 0.905 7.710 1.445 ;
        RECT 5.735 0.735 7.710 0.905 ;
        RECT 5.735 0.725 7.055 0.735 ;
        RECT 5.735 0.255 6.115 0.725 ;
        RECT 6.675 0.255 7.055 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.820 2.805 ;
        RECT 0.145 1.455 0.395 2.635 ;
        RECT 0.615 1.955 0.865 2.465 ;
        RECT 1.085 2.125 1.335 2.635 ;
        RECT 1.555 2.295 2.745 2.465 ;
        RECT 1.555 2.125 1.805 2.295 ;
        RECT 2.495 2.125 2.745 2.295 ;
        RECT 2.965 2.125 3.725 2.635 ;
        RECT 3.945 2.295 5.135 2.465 ;
        RECT 3.945 2.125 4.195 2.295 ;
        RECT 4.885 2.125 5.135 2.295 ;
        RECT 5.355 2.125 5.605 2.635 ;
        RECT 6.295 2.125 6.545 2.635 ;
        RECT 0.615 1.785 5.645 1.955 ;
        RECT 7.235 1.795 7.485 2.635 ;
        RECT 0.085 0.475 0.345 0.895 ;
        RECT 0.615 0.865 0.895 1.785 ;
        RECT 5.475 1.615 5.645 1.785 ;
        RECT 5.475 1.445 5.925 1.615 ;
        RECT 5.705 1.275 5.925 1.445 ;
        RECT 5.705 1.075 7.055 1.275 ;
        RECT 0.515 0.645 0.895 0.865 ;
        RECT 1.115 0.475 1.285 0.905 ;
        RECT 1.455 0.725 5.175 0.905 ;
        RECT 1.455 0.645 4.235 0.725 ;
        RECT 0.085 0.255 3.255 0.475 ;
        RECT 3.435 0.085 3.765 0.465 ;
        RECT 3.985 0.255 4.235 0.645 ;
        RECT 4.455 0.085 4.625 0.555 ;
        RECT 4.795 0.255 5.175 0.725 ;
        RECT 5.395 0.085 5.565 0.905 ;
        RECT 6.335 0.085 6.505 0.555 ;
        RECT 7.275 0.085 7.530 0.565 ;
        RECT 0.000 -0.085 7.820 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o221a_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__o221ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o221ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 3.065 1.075 3.575 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.855 1.615 3.125 2.405 ;
        RECT 2.635 1.445 3.125 1.615 ;
        RECT 2.635 1.245 2.895 1.445 ;
        RECT 2.505 1.075 2.895 1.245 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.015 0.995 1.595 1.325 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 0.995 2.325 1.325 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.465 1.325 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.655 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.974500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.705 0.365 2.465 ;
        RECT 1.900 2.180 2.505 2.465 ;
        RECT 1.900 1.705 2.465 2.180 ;
        RECT 0.085 1.495 2.465 1.705 ;
        RECT 0.675 0.825 0.845 1.495 ;
        RECT 0.085 0.645 0.845 0.825 ;
        RECT 0.085 0.365 0.345 0.645 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.600 1.875 1.580 2.635 ;
        RECT 3.315 1.455 3.575 2.635 ;
        RECT 2.445 0.825 3.575 0.865 ;
        RECT 1.250 0.695 3.575 0.825 ;
        RECT 1.250 0.645 2.560 0.695 ;
        RECT 0.515 0.305 2.065 0.475 ;
        RECT 2.285 0.280 2.560 0.645 ;
        RECT 2.845 0.085 3.015 0.525 ;
        RECT 3.185 0.280 3.575 0.695 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o221ai_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__o221ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o221ai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 3.730 1.445 5.265 1.615 ;
        RECT 3.730 1.075 4.110 1.445 ;
        RECT 5.095 1.275 5.265 1.445 ;
        RECT 5.095 1.075 5.835 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 4.280 1.075 4.875 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 1.120 1.445 3.560 1.615 ;
        RECT 1.120 1.075 2.185 1.445 ;
        RECT 3.180 1.075 3.560 1.445 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 2.355 1.075 3.010 1.275 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.435 1.275 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.105 5.820 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.078000 ;
    PORT
      LAYER li1 ;
        RECT 0.610 1.955 0.860 2.465 ;
        RECT 2.540 1.955 2.790 2.125 ;
        RECT 4.500 1.955 4.750 2.125 ;
        RECT 0.610 1.785 4.750 1.955 ;
        RECT 0.610 1.445 0.900 1.785 ;
        RECT 0.655 0.865 0.900 1.445 ;
        RECT 0.520 0.645 0.900 0.865 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.140 1.455 0.390 2.635 ;
        RECT 1.080 2.125 1.850 2.635 ;
        RECT 2.070 2.295 3.260 2.465 ;
        RECT 2.070 2.125 2.320 2.295 ;
        RECT 3.010 2.125 3.260 2.295 ;
        RECT 3.480 2.125 3.810 2.635 ;
        RECT 4.030 2.295 5.220 2.465 ;
        RECT 4.030 2.125 4.280 2.295 ;
        RECT 4.970 1.785 5.220 2.295 ;
        RECT 5.485 1.455 5.690 2.635 ;
        RECT 0.100 0.475 0.350 0.895 ;
        RECT 1.120 0.645 3.300 0.905 ;
        RECT 3.520 0.735 5.730 0.905 ;
        RECT 1.120 0.475 1.370 0.645 ;
        RECT 3.520 0.475 3.850 0.735 ;
        RECT 4.410 0.725 5.730 0.735 ;
        RECT 0.100 0.255 1.370 0.475 ;
        RECT 1.560 0.255 3.850 0.475 ;
        RECT 4.070 0.085 4.240 0.555 ;
        RECT 4.410 0.255 4.790 0.725 ;
        RECT 5.010 0.085 5.180 0.555 ;
        RECT 5.350 0.255 5.730 0.725 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o221ai_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__o221ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o221ai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.580 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 6.565 1.445 9.320 1.615 ;
        RECT 6.565 1.075 6.945 1.445 ;
        RECT 9.005 1.275 9.320 1.445 ;
        RECT 9.005 1.075 10.135 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 7.125 1.075 8.735 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 4.735 1.445 6.395 1.615 ;
        RECT 4.735 1.275 4.925 1.445 ;
        RECT 2.560 1.075 4.925 1.275 ;
        RECT 6.015 1.075 6.395 1.445 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 5.095 0.995 5.835 1.275 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 1.900 1.275 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.580 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 10.535 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.770 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.580 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.156000 ;
    PORT
      LAYER li1 ;
        RECT 0.625 1.615 0.875 2.465 ;
        RECT 1.565 1.955 1.815 2.465 ;
        RECT 1.565 1.615 2.325 1.955 ;
        RECT 4.345 1.785 8.565 2.005 ;
        RECT 4.345 1.615 4.565 1.785 ;
        RECT 0.625 1.445 4.565 1.615 ;
        RECT 2.120 0.865 2.325 1.445 ;
        RECT 0.535 0.645 2.325 0.865 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.580 2.805 ;
        RECT 0.155 1.485 0.405 2.635 ;
        RECT 1.095 1.825 1.345 2.635 ;
        RECT 2.035 2.125 2.805 2.635 ;
        RECT 3.025 1.955 3.275 2.465 ;
        RECT 3.495 2.125 3.745 2.635 ;
        RECT 3.965 2.265 6.135 2.465 ;
        RECT 3.965 1.955 4.175 2.265 ;
        RECT 6.355 2.175 6.605 2.635 ;
        RECT 6.775 2.265 8.995 2.465 ;
        RECT 3.025 1.785 4.175 1.955 ;
        RECT 8.785 1.955 8.995 2.265 ;
        RECT 9.215 2.125 9.465 2.635 ;
        RECT 9.685 1.955 9.935 2.465 ;
        RECT 8.785 1.785 9.935 1.955 ;
        RECT 9.685 1.445 9.935 1.785 ;
        RECT 10.155 1.445 10.405 2.635 ;
        RECT 0.115 0.475 0.365 0.895 ;
        RECT 6.015 0.820 10.445 0.905 ;
        RECT 2.515 0.735 10.445 0.820 ;
        RECT 2.515 0.645 6.685 0.735 ;
        RECT 0.115 0.255 6.135 0.475 ;
        RECT 6.355 0.255 6.685 0.645 ;
        RECT 7.245 0.725 8.565 0.735 ;
        RECT 6.905 0.085 7.075 0.555 ;
        RECT 7.245 0.255 7.625 0.725 ;
        RECT 7.845 0.085 8.015 0.555 ;
        RECT 8.185 0.255 8.565 0.725 ;
        RECT 9.125 0.725 10.445 0.735 ;
        RECT 8.785 0.085 8.955 0.555 ;
        RECT 9.125 0.255 9.505 0.725 ;
        RECT 9.725 0.085 9.895 0.555 ;
        RECT 10.065 0.255 10.445 0.725 ;
        RECT 0.000 -0.085 10.580 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o221ai_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__or2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__or2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.950 0.765 1.285 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.440 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.005 0.785 1.985 1.015 ;
        RECT 0.010 0.105 1.985 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.551500 ;
    PORT
      LAYER li1 ;
        RECT 1.645 1.845 2.215 2.465 ;
        RECT 1.915 0.825 2.215 1.845 ;
        RECT 1.515 0.255 2.215 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.120 1.665 0.510 1.840 ;
        RECT 1.095 1.835 1.425 2.635 ;
        RECT 0.120 1.495 1.745 1.665 ;
        RECT 0.610 0.595 0.780 1.495 ;
        RECT 1.525 0.995 1.745 1.495 ;
        RECT 0.110 0.085 0.350 0.595 ;
        RECT 0.610 0.265 0.850 0.595 ;
        RECT 1.130 0.085 1.345 0.595 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or2_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__or2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__or2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.915 0.765 1.375 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.765 0.345 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.010 0.785 2.480 1.015 ;
        RECT 0.005 0.105 2.480 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.530500 ;
    PORT
      LAYER li1 ;
        RECT 1.540 2.005 1.920 2.465 ;
        RECT 1.540 1.835 2.415 2.005 ;
        RECT 1.935 0.825 2.415 1.835 ;
        RECT 1.670 0.655 2.415 0.825 ;
        RECT 1.670 0.385 1.840 0.655 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.155 1.665 0.515 1.840 ;
        RECT 1.200 1.835 1.370 2.635 ;
        RECT 2.140 2.175 2.310 2.635 ;
        RECT 0.155 1.495 1.765 1.665 ;
        RECT 0.515 0.595 0.745 1.495 ;
        RECT 1.545 0.995 1.765 1.495 ;
        RECT 0.105 0.085 0.345 0.595 ;
        RECT 0.515 0.255 0.855 0.595 ;
        RECT 1.135 0.085 1.450 0.595 ;
        RECT 2.010 0.085 2.390 0.485 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or2_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__or2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__or2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.915 0.995 1.340 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.765 0.345 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.420 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.028500 ;
    PORT
      LAYER li1 ;
        RECT 1.590 2.005 1.970 2.465 ;
        RECT 2.530 2.005 2.910 2.465 ;
        RECT 1.590 1.835 2.910 2.005 ;
        RECT 2.530 1.665 2.910 1.835 ;
        RECT 2.530 1.495 3.170 1.665 ;
        RECT 2.825 0.905 3.170 1.495 ;
        RECT 1.590 0.735 3.170 0.905 ;
        RECT 1.590 0.265 1.970 0.735 ;
        RECT 2.530 0.265 2.910 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.155 1.665 0.515 2.465 ;
        RECT 1.160 1.835 1.330 2.635 ;
        RECT 2.140 2.175 2.310 2.635 ;
        RECT 3.080 1.835 3.250 2.635 ;
        RECT 0.155 1.495 1.765 1.665 ;
        RECT 0.515 0.825 0.745 1.495 ;
        RECT 1.510 1.245 1.765 1.495 ;
        RECT 1.510 1.075 2.620 1.245 ;
        RECT 0.105 0.085 0.345 0.595 ;
        RECT 0.515 0.290 0.895 0.825 ;
        RECT 1.160 0.085 1.330 0.825 ;
        RECT 2.140 0.085 2.310 0.565 ;
        RECT 3.080 0.085 3.250 0.565 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or2_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__or2_6
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__or2_6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.415 1.075 1.085 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 1.355 1.075 2.025 1.275 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.765 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.396500 ;
    PORT
      LAYER li1 ;
        RECT 2.985 1.665 3.315 2.465 ;
        RECT 3.925 1.665 4.255 2.465 ;
        RECT 4.865 1.665 5.195 2.465 ;
        RECT 2.985 1.495 5.415 1.665 ;
        RECT 5.015 0.905 5.415 1.495 ;
        RECT 2.985 0.725 5.415 0.905 ;
        RECT 2.985 0.255 3.285 0.725 ;
        RECT 3.955 0.255 4.225 0.725 ;
        RECT 4.895 0.255 5.165 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.090 1.665 0.415 2.465 ;
        RECT 0.585 1.835 0.915 2.635 ;
        RECT 1.085 2.295 2.325 2.465 ;
        RECT 1.085 1.665 1.355 2.295 ;
        RECT 0.090 1.455 1.355 1.665 ;
        RECT 1.525 1.665 1.855 2.125 ;
        RECT 2.025 1.835 2.325 2.295 ;
        RECT 1.525 1.445 2.375 1.665 ;
        RECT 2.545 1.495 2.815 2.635 ;
        RECT 3.485 1.835 3.755 2.635 ;
        RECT 4.425 1.835 4.695 2.635 ;
        RECT 5.365 1.835 5.635 2.635 ;
        RECT 2.195 1.275 2.375 1.445 ;
        RECT 2.195 1.075 4.845 1.275 ;
        RECT 2.195 0.905 2.375 1.075 ;
        RECT 0.145 0.085 0.415 0.905 ;
        RECT 0.585 0.735 2.375 0.905 ;
        RECT 0.585 0.725 1.855 0.735 ;
        RECT 0.585 0.255 0.915 0.725 ;
        RECT 1.085 0.085 1.355 0.555 ;
        RECT 1.525 0.255 1.855 0.725 ;
        RECT 2.545 0.555 2.815 0.905 ;
        RECT 2.025 0.085 2.815 0.555 ;
        RECT 3.455 0.085 3.785 0.555 ;
        RECT 4.395 0.085 4.725 0.555 ;
        RECT 5.335 0.085 5.665 0.555 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or2_6

#--------EOF---------

MACRO sky130_fd_sc_hdll__or2_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__or2_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.900 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.415 1.075 1.085 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 1.355 1.075 2.025 1.275 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.900 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 6.705 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.090 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.900 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.862000 ;
    PORT
      LAYER li1 ;
        RECT 2.985 1.665 3.315 2.465 ;
        RECT 3.925 1.665 4.255 2.465 ;
        RECT 4.865 1.665 5.195 2.465 ;
        RECT 5.805 1.665 6.135 2.465 ;
        RECT 2.985 1.495 6.335 1.665 ;
        RECT 5.935 0.905 6.335 1.495 ;
        RECT 2.985 0.725 6.335 0.905 ;
        RECT 2.985 0.255 3.285 0.725 ;
        RECT 3.955 0.255 4.225 0.725 ;
        RECT 4.895 0.255 5.165 0.725 ;
        RECT 5.835 0.255 6.105 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.900 2.805 ;
        RECT 0.090 1.665 0.415 2.465 ;
        RECT 0.585 1.835 0.915 2.635 ;
        RECT 1.085 2.295 2.325 2.465 ;
        RECT 1.085 1.665 1.355 2.295 ;
        RECT 0.090 1.455 1.355 1.665 ;
        RECT 1.525 1.665 1.855 2.125 ;
        RECT 2.025 1.835 2.325 2.295 ;
        RECT 1.525 1.445 2.375 1.665 ;
        RECT 2.545 1.495 2.815 2.635 ;
        RECT 3.485 1.835 3.755 2.635 ;
        RECT 4.425 1.835 4.695 2.635 ;
        RECT 5.365 1.835 5.635 2.635 ;
        RECT 6.305 1.835 6.575 2.635 ;
        RECT 2.195 1.275 2.375 1.445 ;
        RECT 2.195 1.075 5.525 1.275 ;
        RECT 2.195 0.905 2.375 1.075 ;
        RECT 0.145 0.085 0.415 0.905 ;
        RECT 0.585 0.735 2.375 0.905 ;
        RECT 0.585 0.725 1.855 0.735 ;
        RECT 0.585 0.255 0.915 0.725 ;
        RECT 1.085 0.085 1.355 0.555 ;
        RECT 1.525 0.255 1.855 0.725 ;
        RECT 2.545 0.555 2.815 0.905 ;
        RECT 2.025 0.085 2.815 0.555 ;
        RECT 3.455 0.085 3.785 0.555 ;
        RECT 4.395 0.085 4.725 0.555 ;
        RECT 5.335 0.085 5.665 0.555 ;
        RECT 6.275 0.085 6.605 0.555 ;
        RECT 0.000 -0.085 6.900 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or2_8

#--------EOF---------

MACRO sky130_fd_sc_hdll__or2b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__or2b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.540 2.085 1.835 2.415 ;
    END
  END A
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 0.425 1.325 ;
    END
  END B_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.960 0.815 2.955 1.015 ;
        RECT 0.005 0.135 2.955 0.815 ;
        RECT 0.150 -0.085 0.320 0.135 ;
        RECT 1.960 0.105 2.955 0.135 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.455500 ;
    PORT
      LAYER li1 ;
        RECT 2.605 1.495 3.090 2.465 ;
        RECT 2.705 0.760 3.090 1.495 ;
        RECT 2.605 0.415 3.090 0.760 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.090 1.495 0.345 2.635 ;
        RECT 0.645 1.325 0.815 1.885 ;
        RECT 1.040 1.665 1.460 1.915 ;
        RECT 2.065 1.835 2.345 2.635 ;
        RECT 1.040 1.495 2.385 1.665 ;
        RECT 2.215 1.325 2.385 1.495 ;
        RECT 0.645 0.995 1.385 1.325 ;
        RECT 2.215 0.995 2.445 1.325 ;
        RECT 0.645 0.905 0.895 0.995 ;
        RECT 0.110 0.735 0.895 0.905 ;
        RECT 2.215 0.825 2.385 0.995 ;
        RECT 0.110 0.265 0.420 0.735 ;
        RECT 1.595 0.655 2.385 0.825 ;
        RECT 0.640 0.085 1.375 0.565 ;
        RECT 1.595 0.305 1.765 0.655 ;
        RECT 1.935 0.085 2.365 0.485 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or2b_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__or2b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__or2b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.540 2.085 1.830 2.415 ;
    END
  END A
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.425 1.325 ;
    END
  END B_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.955 0.815 3.625 1.015 ;
        RECT 0.005 0.135 3.625 0.815 ;
        RECT 0.145 -0.085 0.315 0.135 ;
        RECT 1.955 0.105 3.625 0.135 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.811500 ;
    PORT
      LAYER li1 ;
        RECT 2.790 0.415 3.110 2.465 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.085 1.495 0.345 2.635 ;
        RECT 0.645 1.325 0.815 1.885 ;
        RECT 1.035 1.665 1.455 1.915 ;
        RECT 2.060 1.835 2.340 2.635 ;
        RECT 1.035 1.495 2.440 1.665 ;
        RECT 0.645 0.995 1.380 1.325 ;
        RECT 0.645 0.905 0.890 0.995 ;
        RECT 0.105 0.735 0.890 0.905 ;
        RECT 2.270 0.825 2.440 1.495 ;
        RECT 3.285 1.460 3.520 2.635 ;
        RECT 0.105 0.265 0.420 0.735 ;
        RECT 1.590 0.655 2.440 0.825 ;
        RECT 0.640 0.085 1.370 0.565 ;
        RECT 1.590 0.305 1.760 0.655 ;
        RECT 2.030 0.085 2.360 0.485 ;
        RECT 3.285 0.085 3.520 0.925 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or2b_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__or2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__or2b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.730 1.075 2.470 1.275 ;
    END
  END A
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 0.425 1.955 ;
    END
  END B_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.830 0.815 4.425 1.015 ;
        RECT 0.005 0.135 4.425 0.815 ;
        RECT 0.145 0.105 4.425 0.135 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.028500 ;
    PORT
      LAYER li1 ;
        RECT 2.565 1.955 2.815 2.465 ;
        RECT 3.505 1.955 3.755 2.465 ;
        RECT 2.565 1.785 3.755 1.955 ;
        RECT 3.080 1.615 3.755 1.785 ;
        RECT 3.080 1.445 4.490 1.615 ;
        RECT 4.105 0.905 4.490 1.445 ;
        RECT 2.475 0.735 4.490 0.905 ;
        RECT 2.475 0.290 2.855 0.735 ;
        RECT 3.415 0.290 3.795 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.090 2.125 0.345 2.635 ;
        RECT 0.645 1.325 0.815 2.465 ;
        RECT 1.040 1.615 1.560 2.465 ;
        RECT 2.065 1.835 2.345 2.635 ;
        RECT 3.035 2.135 3.285 2.635 ;
        RECT 3.975 1.795 4.225 2.635 ;
        RECT 1.040 1.495 2.860 1.615 ;
        RECT 1.340 1.445 2.860 1.495 ;
        RECT 0.645 0.995 1.170 1.325 ;
        RECT 0.645 0.905 0.895 0.995 ;
        RECT 0.110 0.735 0.895 0.905 ;
        RECT 1.340 0.905 1.560 1.445 ;
        RECT 2.690 1.245 2.860 1.445 ;
        RECT 2.690 1.075 3.800 1.245 ;
        RECT 1.340 0.735 1.845 0.905 ;
        RECT 0.110 0.265 0.420 0.735 ;
        RECT 0.640 0.085 1.295 0.565 ;
        RECT 1.465 0.305 1.845 0.735 ;
        RECT 2.130 0.085 2.305 0.905 ;
        RECT 3.075 0.085 3.245 0.550 ;
        RECT 4.015 0.085 4.185 0.550 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or2b_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__or3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__or3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.325 0.845 1.615 ;
        RECT 0.605 0.995 1.490 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.085 2.125 1.375 2.415 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.430 1.325 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.490 0.815 2.700 1.015 ;
        RECT 0.015 0.135 2.700 0.815 ;
        RECT 0.140 -0.085 0.310 0.135 ;
        RECT 1.490 0.105 2.700 0.135 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.810250 ;
    PORT
      LAYER li1 ;
        RECT 2.340 1.495 2.615 2.465 ;
        RECT 2.445 0.760 2.615 1.495 ;
        RECT 2.340 0.415 2.615 0.760 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.105 1.785 1.375 1.955 ;
        RECT 1.595 1.835 1.875 2.635 ;
        RECT 0.105 1.495 0.430 1.785 ;
        RECT 1.205 1.665 1.375 1.785 ;
        RECT 1.205 1.495 1.975 1.665 ;
        RECT 1.805 0.825 1.975 1.495 ;
        RECT 0.100 0.655 1.975 0.825 ;
        RECT 0.100 0.305 0.355 0.655 ;
        RECT 0.525 0.085 0.905 0.485 ;
        RECT 1.125 0.305 1.295 0.655 ;
        RECT 1.465 0.085 1.895 0.485 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or3_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__or3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__or3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.555 1.325 0.880 1.615 ;
        RECT 0.555 0.995 1.580 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.085 2.125 1.380 2.415 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.385 1.325 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.495 0.815 3.165 1.015 ;
        RECT 0.020 0.135 3.165 0.815 ;
        RECT 0.145 -0.085 0.315 0.135 ;
        RECT 1.495 0.105 3.165 0.135 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.530500 ;
    PORT
      LAYER li1 ;
        RECT 2.330 1.495 2.655 2.465 ;
        RECT 2.470 0.760 2.655 1.495 ;
        RECT 2.330 0.415 2.655 0.760 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.105 1.785 1.370 1.955 ;
        RECT 1.600 1.835 2.070 2.635 ;
        RECT 0.105 1.495 0.385 1.785 ;
        RECT 1.200 1.665 1.370 1.785 ;
        RECT 1.200 1.495 2.110 1.665 ;
        RECT 1.890 1.325 2.110 1.495 ;
        RECT 2.825 1.430 3.115 2.635 ;
        RECT 1.890 0.995 2.300 1.325 ;
        RECT 1.890 0.825 2.110 0.995 ;
        RECT 0.105 0.655 2.110 0.825 ;
        RECT 0.105 0.305 0.360 0.655 ;
        RECT 0.530 0.085 0.910 0.485 ;
        RECT 1.130 0.305 1.300 0.655 ;
        RECT 1.470 0.085 2.090 0.485 ;
        RECT 2.825 0.085 3.115 0.915 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or3_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__or3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__or3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.325 1.075 1.850 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.595 1.325 0.830 2.050 ;
        RECT 0.595 1.075 1.155 1.325 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.425 1.325 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.390 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.996000 ;
    PORT
      LAYER li1 ;
        RECT 2.545 1.615 2.795 2.465 ;
        RECT 3.485 1.615 3.735 2.465 ;
        RECT 2.545 1.445 4.455 1.615 ;
        RECT 4.115 0.905 4.455 1.445 ;
        RECT 2.455 0.735 4.455 0.905 ;
        RECT 2.455 0.265 2.835 0.735 ;
        RECT 3.395 0.265 3.775 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.085 2.295 1.365 2.465 ;
        RECT 0.085 1.495 0.425 2.295 ;
        RECT 1.100 1.665 1.365 2.295 ;
        RECT 1.585 1.835 2.285 2.635 ;
        RECT 3.015 1.795 3.265 2.635 ;
        RECT 3.955 1.795 4.205 2.635 ;
        RECT 1.100 1.495 2.240 1.665 ;
        RECT 2.020 1.245 2.240 1.495 ;
        RECT 2.020 1.075 3.945 1.245 ;
        RECT 2.020 0.905 2.240 1.075 ;
        RECT 0.085 0.725 2.240 0.905 ;
        RECT 0.085 0.255 0.425 0.725 ;
        RECT 0.645 0.085 0.815 0.555 ;
        RECT 0.985 0.255 1.365 0.725 ;
        RECT 1.585 0.085 2.285 0.555 ;
        RECT 3.055 0.085 3.225 0.555 ;
        RECT 3.995 0.085 4.165 0.555 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or3_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__or3b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__or3b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.525 1.325 1.770 1.615 ;
        RECT 1.525 0.995 2.465 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.635 2.125 2.350 2.455 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 0.425 1.325 ;
    END
  END C_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.815 0.985 1.015 ;
        RECT 2.470 0.815 3.465 1.015 ;
        RECT 0.005 0.335 3.465 0.815 ;
        RECT 0.145 0.135 3.465 0.335 ;
        RECT 0.145 -0.085 0.315 0.135 ;
        RECT 2.470 0.105 3.465 0.135 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.463750 ;
    PORT
      LAYER li1 ;
        RECT 3.110 1.495 3.535 2.465 ;
        RECT 3.215 0.760 3.535 1.495 ;
        RECT 3.110 0.415 3.535 0.760 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.085 1.495 0.345 2.635 ;
        RECT 0.645 1.325 0.815 1.885 ;
        RECT 1.075 1.785 2.350 1.955 ;
        RECT 2.570 1.835 2.850 2.635 ;
        RECT 1.075 1.495 1.335 1.785 ;
        RECT 2.180 1.665 2.350 1.785 ;
        RECT 2.180 1.495 2.890 1.665 ;
        RECT 2.720 1.325 2.890 1.495 ;
        RECT 0.645 0.995 1.270 1.325 ;
        RECT 2.720 0.995 2.995 1.325 ;
        RECT 0.645 0.905 0.895 0.995 ;
        RECT 0.085 0.085 0.345 0.905 ;
        RECT 0.515 0.485 0.895 0.905 ;
        RECT 2.720 0.825 2.890 0.995 ;
        RECT 1.075 0.655 2.890 0.825 ;
        RECT 1.075 0.255 1.335 0.655 ;
        RECT 1.505 0.085 1.885 0.485 ;
        RECT 2.105 0.305 2.275 0.655 ;
        RECT 2.445 0.085 2.870 0.485 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or3b_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__or3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__or3b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.955 1.075 2.540 1.615 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 2.195 2.125 3.545 2.365 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.425 1.640 ;
    END
  END C_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.540 0.815 2.135 1.015 ;
        RECT 0.540 0.785 3.580 0.815 ;
        RECT 0.005 0.135 3.580 0.785 ;
        RECT 0.005 0.105 2.190 0.135 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.741250 ;
    PORT
      LAYER li1 ;
        RECT 0.985 1.495 1.430 1.700 ;
        RECT 0.985 0.595 1.235 1.495 ;
        RECT 0.985 0.265 1.385 0.595 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.085 2.040 0.345 2.220 ;
        RECT 0.600 2.210 0.960 2.635 ;
        RECT 1.685 2.210 2.015 2.635 ;
        RECT 0.085 1.955 1.980 2.040 ;
        RECT 0.085 1.870 3.020 1.955 ;
        RECT 0.085 1.810 0.815 1.870 ;
        RECT 0.645 0.905 0.815 1.810 ;
        RECT 1.810 1.785 3.020 1.870 ;
        RECT 2.850 1.325 3.020 1.785 ;
        RECT 3.240 1.495 3.545 1.925 ;
        RECT 0.085 0.735 0.815 0.905 ;
        RECT 1.485 0.905 1.655 1.325 ;
        RECT 2.850 0.995 3.200 1.325 ;
        RECT 1.485 0.825 2.535 0.905 ;
        RECT 3.375 0.825 3.545 1.495 ;
        RECT 1.485 0.735 3.545 0.825 ;
        RECT 0.085 0.290 0.345 0.735 ;
        RECT 2.365 0.655 3.545 0.735 ;
        RECT 0.645 0.085 0.815 0.565 ;
        RECT 1.865 0.085 2.035 0.565 ;
        RECT 2.365 0.305 2.535 0.655 ;
        RECT 2.740 0.085 3.070 0.485 ;
        RECT 3.240 0.305 3.545 0.655 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or3b_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__or3b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__or3b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.800 0.995 3.110 1.700 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 3.330 0.995 3.570 1.700 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.425 1.640 ;
    END
  END C_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.540 0.785 4.400 1.015 ;
        RECT 0.005 0.105 4.400 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.028500 ;
    PORT
      LAYER li1 ;
        RECT 1.010 1.415 2.420 1.700 ;
        RECT 1.010 0.905 1.270 1.415 ;
        RECT 1.010 0.735 2.240 0.905 ;
        RECT 1.010 0.285 1.430 0.735 ;
        RECT 2.005 0.255 2.240 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.085 2.040 0.345 2.220 ;
        RECT 0.600 2.210 0.960 2.635 ;
        RECT 1.520 2.210 1.900 2.635 ;
        RECT 2.455 2.210 2.845 2.635 ;
        RECT 3.870 2.210 4.455 2.425 ;
        RECT 0.085 1.870 4.030 2.040 ;
        RECT 0.085 1.810 0.815 1.870 ;
        RECT 0.645 0.905 0.815 1.810 ;
        RECT 1.440 1.075 2.615 1.245 ;
        RECT 0.085 0.735 0.815 0.905 ;
        RECT 2.445 0.825 2.615 1.075 ;
        RECT 3.860 0.995 4.030 1.870 ;
        RECT 4.250 0.825 4.455 2.210 ;
        RECT 0.085 0.290 0.345 0.735 ;
        RECT 2.445 0.655 4.455 0.825 ;
        RECT 0.670 0.085 0.840 0.565 ;
        RECT 1.650 0.085 1.820 0.565 ;
        RECT 2.460 0.085 2.840 0.485 ;
        RECT 3.400 0.085 3.840 0.485 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or3b_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__or4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__or4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.525 0.995 2.095 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.090 2.125 1.895 2.415 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.660 0.995 1.355 1.615 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.755 0.440 1.325 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.010 0.815 3.155 1.015 ;
        RECT 0.005 0.135 3.155 0.815 ;
        RECT 0.150 -0.085 0.320 0.135 ;
        RECT 2.010 0.105 3.155 0.135 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.703000 ;
    PORT
      LAYER li1 ;
        RECT 2.805 1.495 3.075 2.465 ;
        RECT 2.905 0.760 3.075 1.495 ;
        RECT 2.805 0.415 3.075 0.760 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.090 1.785 1.830 1.955 ;
        RECT 2.115 1.835 2.395 2.635 ;
        RECT 0.090 1.495 0.410 1.785 ;
        RECT 1.660 1.665 1.830 1.785 ;
        RECT 1.660 1.495 2.435 1.665 ;
        RECT 2.265 1.325 2.435 1.495 ;
        RECT 2.265 0.995 2.555 1.325 ;
        RECT 2.265 0.825 2.435 0.995 ;
        RECT 0.675 0.655 2.435 0.825 ;
        RECT 0.095 0.085 0.425 0.585 ;
        RECT 0.675 0.305 0.845 0.655 ;
        RECT 1.045 0.085 1.425 0.485 ;
        RECT 1.645 0.305 1.815 0.655 ;
        RECT 1.985 0.085 2.415 0.485 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or4_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__or4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__or4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.475 0.995 2.095 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.085 2.125 1.895 2.415 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.995 1.305 1.615 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.755 0.435 1.325 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.010 0.815 3.675 1.015 ;
        RECT 0.005 0.135 3.675 0.815 ;
        RECT 0.150 -0.085 0.320 0.135 ;
        RECT 2.010 0.105 3.675 0.135 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.802750 ;
    PORT
      LAYER li1 ;
        RECT 2.820 1.495 3.125 2.465 ;
        RECT 2.890 0.760 3.125 1.495 ;
        RECT 2.820 0.415 3.125 0.760 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.085 1.785 1.830 1.955 ;
        RECT 2.115 1.835 2.395 2.635 ;
        RECT 0.085 1.495 0.410 1.785 ;
        RECT 1.660 1.665 1.830 1.785 ;
        RECT 1.660 1.495 2.435 1.665 ;
        RECT 2.265 1.325 2.435 1.495 ;
        RECT 3.315 1.455 3.535 2.635 ;
        RECT 2.265 0.995 2.700 1.325 ;
        RECT 2.265 0.825 2.435 0.995 ;
        RECT 0.675 0.655 2.435 0.825 ;
        RECT 0.090 0.085 0.425 0.585 ;
        RECT 0.675 0.305 0.845 0.655 ;
        RECT 1.045 0.085 1.425 0.485 ;
        RECT 1.645 0.305 1.815 0.655 ;
        RECT 1.985 0.085 2.415 0.485 ;
        RECT 3.315 0.085 3.535 1.000 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or4_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__or4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__or4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.940 1.445 2.475 1.615 ;
        RECT 1.940 0.995 2.210 1.445 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.500 1.785 1.870 2.375 ;
        RECT 1.500 1.450 1.760 1.785 ;
        RECT 1.380 0.995 1.760 1.450 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.930 1.620 1.330 2.375 ;
        RECT 0.930 0.995 1.100 1.620 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.755 0.370 1.325 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.030 0.105 4.535 1.015 ;
        RECT 0.140 -0.085 0.310 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.028500 ;
    PORT
      LAYER li1 ;
        RECT 2.730 1.625 2.980 2.465 ;
        RECT 3.670 1.625 3.920 2.465 ;
        RECT 2.730 1.455 4.485 1.625 ;
        RECT 4.210 0.905 4.485 1.455 ;
        RECT 2.770 0.725 4.485 0.905 ;
        RECT 2.770 0.255 3.020 0.725 ;
        RECT 3.580 0.255 3.960 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.115 1.665 0.450 2.450 ;
        RECT 2.205 1.795 2.455 2.635 ;
        RECT 3.200 1.795 3.450 2.635 ;
        RECT 4.140 1.795 4.390 2.635 ;
        RECT 0.115 1.495 0.760 1.665 ;
        RECT 0.540 0.825 0.760 1.495 ;
        RECT 2.380 1.075 3.990 1.245 ;
        RECT 2.380 0.825 2.550 1.075 ;
        RECT 0.540 0.655 2.550 0.825 ;
        RECT 0.120 0.085 0.370 0.585 ;
        RECT 0.750 0.305 0.920 0.655 ;
        RECT 1.120 0.085 1.500 0.485 ;
        RECT 1.720 0.305 1.890 0.655 ;
        RECT 2.160 0.085 2.540 0.485 ;
        RECT 3.240 0.085 3.410 0.555 ;
        RECT 4.180 0.085 4.350 0.555 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or4_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__or4b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__or4b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 2.630 0.995 3.075 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.660 2.125 2.860 2.415 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.620 0.995 2.410 1.615 ;
    END
  END C
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.755 0.425 1.325 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.975 0.815 3.975 1.015 ;
        RECT 0.005 0.135 3.975 0.815 ;
        RECT 0.150 -0.085 0.320 0.135 ;
        RECT 2.975 0.105 3.975 0.135 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.463750 ;
    PORT
      LAYER li1 ;
        RECT 3.620 1.495 3.995 2.465 ;
        RECT 3.725 0.760 3.995 1.495 ;
        RECT 3.620 0.415 3.995 0.760 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.085 1.560 0.425 2.635 ;
        RECT 0.645 1.325 0.885 1.920 ;
        RECT 1.080 1.785 2.860 1.955 ;
        RECT 3.080 1.835 3.360 2.635 ;
        RECT 1.080 1.495 1.400 1.785 ;
        RECT 2.690 1.665 2.860 1.785 ;
        RECT 2.690 1.495 3.415 1.665 ;
        RECT 3.245 1.325 3.415 1.495 ;
        RECT 0.645 0.995 1.300 1.325 ;
        RECT 3.245 0.995 3.505 1.325 ;
        RECT 0.085 0.085 0.425 0.585 ;
        RECT 0.645 0.305 0.890 0.995 ;
        RECT 3.245 0.825 3.415 0.995 ;
        RECT 1.665 0.655 3.415 0.825 ;
        RECT 1.085 0.085 1.415 0.585 ;
        RECT 1.665 0.305 1.835 0.655 ;
        RECT 2.010 0.085 2.390 0.485 ;
        RECT 2.610 0.305 2.780 0.655 ;
        RECT 2.950 0.085 3.380 0.485 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or4b_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__or4b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__or4b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.905 1.075 2.520 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 2.185 2.125 2.920 2.415 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 2.800 1.075 3.900 1.275 ;
    END
  END C
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.425 1.435 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.540 0.785 1.990 1.015 ;
        RECT 0.005 0.105 3.995 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.498000 ;
    PORT
      LAYER li1 ;
        RECT 1.020 1.495 1.350 1.825 ;
        RECT 1.020 0.790 1.235 1.495 ;
        RECT 1.020 0.260 1.350 0.790 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.515 2.335 0.895 2.635 ;
        RECT 1.630 2.335 1.965 2.635 ;
        RECT 3.160 2.215 3.695 2.385 ;
        RECT 0.510 1.995 1.865 2.165 ;
        RECT 0.510 1.890 0.815 1.995 ;
        RECT 0.085 1.605 0.815 1.890 ;
        RECT 1.540 1.955 1.865 1.995 ;
        RECT 3.160 1.955 3.330 2.215 ;
        RECT 1.540 1.785 3.330 1.955 ;
        RECT 3.525 1.615 3.910 1.780 ;
        RECT 0.645 0.905 0.815 1.605 ;
        RECT 1.520 1.445 3.910 1.615 ;
        RECT 1.520 1.325 1.735 1.445 ;
        RECT 1.405 0.960 1.735 1.325 ;
        RECT 0.085 0.735 0.815 0.905 ;
        RECT 1.565 0.870 1.735 0.960 ;
        RECT 0.085 0.325 0.350 0.735 ;
        RECT 1.565 0.700 3.305 0.870 ;
        RECT 0.680 0.085 0.850 0.565 ;
        RECT 1.535 0.085 1.965 0.485 ;
        RECT 2.185 0.270 2.355 0.700 ;
        RECT 2.585 0.085 2.915 0.485 ;
        RECT 3.135 0.270 3.305 0.700 ;
        RECT 3.525 0.085 3.905 0.585 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or4b_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__or4b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__or4b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.875 1.445 3.440 1.615 ;
        RECT 2.875 0.995 3.175 1.445 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.375 0.995 2.705 2.375 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 1.895 0.995 2.185 2.375 ;
    END
  END C
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.995 0.445 1.955 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.335 5.500 1.015 ;
        RECT 0.145 0.105 5.500 0.335 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.028500 ;
    PORT
      LAYER li1 ;
        RECT 3.695 1.625 3.945 2.465 ;
        RECT 4.635 1.625 4.885 2.465 ;
        RECT 3.695 1.455 5.415 1.625 ;
        RECT 5.175 0.905 5.415 1.455 ;
        RECT 3.735 0.725 5.415 0.905 ;
        RECT 3.735 0.255 3.985 0.725 ;
        RECT 4.545 0.255 4.925 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.085 2.135 0.365 2.635 ;
        RECT 0.645 1.325 0.835 2.455 ;
        RECT 1.085 1.745 1.415 2.450 ;
        RECT 3.170 1.795 3.420 2.635 ;
        RECT 4.165 1.795 4.415 2.635 ;
        RECT 5.105 1.795 5.355 2.635 ;
        RECT 1.085 1.575 1.725 1.745 ;
        RECT 0.645 0.995 1.265 1.325 ;
        RECT 0.085 0.085 0.345 0.825 ;
        RECT 0.645 0.435 0.835 0.995 ;
        RECT 1.505 0.825 1.725 1.575 ;
        RECT 3.345 1.075 4.955 1.245 ;
        RECT 3.345 0.825 3.515 1.075 ;
        RECT 1.505 0.655 3.515 0.825 ;
        RECT 1.085 0.085 1.335 0.585 ;
        RECT 1.715 0.305 1.885 0.655 ;
        RECT 2.085 0.085 2.465 0.485 ;
        RECT 2.685 0.305 2.855 0.655 ;
        RECT 3.125 0.085 3.505 0.485 ;
        RECT 4.205 0.085 4.375 0.555 ;
        RECT 5.145 0.085 5.315 0.555 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or4b_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__or4bb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__or4bb_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 2.815 0.995 3.570 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 2.680 2.125 3.370 2.455 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.995 0.810 1.695 ;
    END
  END C_N
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.980 0.995 1.335 1.325 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.040 0.785 1.515 1.015 ;
        RECT 3.485 0.785 4.485 1.015 ;
        RECT 0.040 0.335 4.485 0.785 ;
        RECT 0.145 -0.085 0.315 0.335 ;
        RECT 1.525 0.105 4.485 0.335 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.463750 ;
    PORT
      LAYER li1 ;
        RECT 4.130 1.495 4.455 2.465 ;
        RECT 4.235 0.760 4.455 1.495 ;
        RECT 4.130 0.415 4.455 0.760 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.085 2.035 0.345 2.455 ;
        RECT 0.515 2.205 0.895 2.635 ;
        RECT 1.610 2.205 2.405 2.375 ;
        RECT 0.085 1.865 2.015 2.035 ;
        RECT 0.085 0.825 0.255 1.865 ;
        RECT 1.040 1.525 1.675 1.695 ;
        RECT 1.505 1.245 1.675 1.525 ;
        RECT 1.845 1.585 2.015 1.865 ;
        RECT 2.235 1.955 2.405 2.205 ;
        RECT 2.235 1.785 3.370 1.955 ;
        RECT 3.590 1.835 3.870 2.635 ;
        RECT 3.200 1.665 3.370 1.785 ;
        RECT 1.845 1.415 2.545 1.585 ;
        RECT 3.200 1.495 3.910 1.665 ;
        RECT 1.505 1.075 2.155 1.245 ;
        RECT 1.505 0.825 1.675 1.075 ;
        RECT 2.375 0.995 2.545 1.415 ;
        RECT 3.740 1.325 3.910 1.495 ;
        RECT 3.740 0.995 4.030 1.325 ;
        RECT 3.740 0.825 3.910 0.995 ;
        RECT 0.085 0.450 0.400 0.825 ;
        RECT 0.705 0.085 0.875 0.825 ;
        RECT 1.175 0.655 1.675 0.825 ;
        RECT 2.165 0.655 3.910 0.825 ;
        RECT 1.175 0.450 1.345 0.655 ;
        RECT 1.570 0.085 1.945 0.485 ;
        RECT 2.165 0.305 2.335 0.655 ;
        RECT 2.520 0.085 2.900 0.485 ;
        RECT 3.120 0.305 3.290 0.655 ;
        RECT 3.460 0.085 3.890 0.485 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or4bb_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__or4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__or4bb_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 2.840 0.995 3.595 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 2.705 2.125 3.395 2.455 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.430 0.995 0.830 1.695 ;
    END
  END C_N
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 1.000 0.995 1.340 1.325 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.045 0.785 1.520 1.015 ;
        RECT 3.510 0.785 4.990 1.015 ;
        RECT 0.045 0.335 4.990 0.785 ;
        RECT 0.150 -0.085 0.320 0.335 ;
        RECT 1.530 0.105 4.990 0.335 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.498000 ;
    PORT
      LAYER li1 ;
        RECT 4.155 1.495 4.455 2.465 ;
        RECT 4.260 0.760 4.455 1.495 ;
        RECT 4.155 0.415 4.455 0.760 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.060 2.805 ;
        RECT 0.085 2.035 0.345 2.455 ;
        RECT 0.515 2.205 0.895 2.635 ;
        RECT 1.635 2.205 2.430 2.375 ;
        RECT 0.085 1.865 2.040 2.035 ;
        RECT 0.085 0.825 0.260 1.865 ;
        RECT 1.045 1.525 1.700 1.695 ;
        RECT 1.510 1.245 1.700 1.525 ;
        RECT 1.870 1.585 2.040 1.865 ;
        RECT 2.260 1.955 2.430 2.205 ;
        RECT 2.260 1.785 3.395 1.955 ;
        RECT 3.615 1.835 3.895 2.635 ;
        RECT 3.225 1.665 3.395 1.785 ;
        RECT 1.870 1.415 2.570 1.585 ;
        RECT 3.225 1.495 3.935 1.665 ;
        RECT 1.510 1.075 1.955 1.245 ;
        RECT 1.510 0.825 1.700 1.075 ;
        RECT 2.400 0.995 2.570 1.415 ;
        RECT 3.765 1.325 3.935 1.495 ;
        RECT 4.650 1.440 4.820 2.635 ;
        RECT 3.765 0.995 4.040 1.325 ;
        RECT 3.765 0.825 3.935 0.995 ;
        RECT 0.085 0.450 0.405 0.825 ;
        RECT 0.710 0.085 0.880 0.825 ;
        RECT 1.180 0.655 1.700 0.825 ;
        RECT 2.190 0.655 3.935 0.825 ;
        RECT 1.180 0.450 1.350 0.655 ;
        RECT 1.595 0.085 1.970 0.485 ;
        RECT 2.190 0.305 2.360 0.655 ;
        RECT 2.545 0.085 2.925 0.485 ;
        RECT 3.145 0.305 3.315 0.655 ;
        RECT 3.485 0.085 3.915 0.485 ;
        RECT 4.650 0.085 4.820 0.915 ;
        RECT 0.000 -0.085 5.060 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or4bb_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__or4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__or4bb_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 3.315 1.400 3.675 1.615 ;
        RECT 3.455 0.995 3.675 1.400 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 2.845 0.995 3.145 2.375 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.435 0.995 0.825 1.695 ;
    END
  END C_N
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 0.995 0.995 1.335 1.325 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.040 0.335 5.975 1.015 ;
        RECT 0.145 -0.085 0.315 0.335 ;
        RECT 1.525 0.105 5.975 0.335 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.285 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.028500 ;
    PORT
      LAYER li1 ;
        RECT 4.185 1.625 4.435 2.465 ;
        RECT 5.125 1.625 5.375 2.465 ;
        RECT 4.185 1.455 5.855 1.625 ;
        RECT 5.625 0.905 5.855 1.455 ;
        RECT 4.225 0.725 5.855 0.905 ;
        RECT 4.225 0.255 4.475 0.725 ;
        RECT 5.035 0.255 5.415 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.095 2.070 0.345 2.455 ;
        RECT 0.515 2.240 0.895 2.635 ;
        RECT 1.225 2.295 2.565 2.465 ;
        RECT 1.225 2.070 1.395 2.295 ;
        RECT 0.095 1.900 1.395 2.070 ;
        RECT 1.610 1.955 2.225 2.125 ;
        RECT 0.095 0.825 0.265 1.900 ;
        RECT 1.040 1.560 1.695 1.730 ;
        RECT 1.505 1.325 1.695 1.560 ;
        RECT 1.505 0.995 1.795 1.325 ;
        RECT 1.505 0.825 1.695 0.995 ;
        RECT 0.095 0.450 0.400 0.825 ;
        RECT 0.705 0.085 0.875 0.825 ;
        RECT 1.175 0.655 1.695 0.825 ;
        RECT 2.035 0.825 2.225 1.955 ;
        RECT 2.395 0.995 2.565 2.295 ;
        RECT 3.660 1.795 3.910 2.635 ;
        RECT 4.655 1.795 4.905 2.635 ;
        RECT 5.595 1.795 5.845 2.635 ;
        RECT 3.845 1.075 5.445 1.245 ;
        RECT 3.845 0.825 4.015 1.075 ;
        RECT 2.035 0.655 4.015 0.825 ;
        RECT 1.175 0.450 1.345 0.655 ;
        RECT 1.615 0.085 1.945 0.480 ;
        RECT 2.245 0.305 2.415 0.655 ;
        RECT 2.585 0.085 2.965 0.485 ;
        RECT 3.185 0.305 3.355 0.655 ;
        RECT 3.615 0.085 3.995 0.485 ;
        RECT 4.695 0.085 4.865 0.555 ;
        RECT 5.635 0.085 5.805 0.555 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or4bb_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__probe_p_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__probe_p_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.832500 ;
    PORT
      LAYER li1 ;
        RECT 0.140 1.075 1.240 1.275 ;
    END
  END A
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.635 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1.250 1.950 4.270 2.160 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.095 1.615 0.425 2.465 ;
        RECT 0.595 1.835 0.865 2.635 ;
        RECT 1.035 1.615 1.365 2.465 ;
        RECT 1.535 1.835 1.805 2.635 ;
        RECT 1.975 1.615 2.305 2.465 ;
        RECT 2.475 1.835 2.745 2.635 ;
        RECT 2.915 1.615 3.245 2.465 ;
        RECT 3.415 1.835 3.685 2.635 ;
        RECT 3.855 1.615 4.185 2.465 ;
        RECT 4.355 1.835 4.625 2.635 ;
        RECT 4.795 1.615 5.125 2.465 ;
        RECT 0.095 1.445 1.595 1.615 ;
        RECT 1.975 1.445 5.125 1.615 ;
        RECT 5.295 1.485 5.595 2.635 ;
        RECT 1.420 1.245 1.595 1.445 ;
        RECT 1.420 1.075 4.045 1.245 ;
        RECT 1.420 0.905 1.595 1.075 ;
        RECT 4.290 0.905 5.125 1.445 ;
        RECT 0.145 0.735 1.595 0.905 ;
        RECT 1.975 0.735 5.125 0.905 ;
        RECT 0.145 0.255 0.445 0.735 ;
        RECT 0.615 0.085 0.895 0.565 ;
        RECT 1.065 0.255 1.335 0.735 ;
        RECT 1.505 0.085 1.805 0.565 ;
        RECT 1.975 0.255 2.305 0.735 ;
        RECT 2.475 0.085 2.745 0.565 ;
        RECT 2.915 0.255 3.245 0.735 ;
        RECT 3.415 0.085 3.685 0.565 ;
        RECT 3.855 0.255 4.185 0.735 ;
        RECT 4.355 0.085 4.625 0.565 ;
        RECT 4.795 0.255 5.125 0.735 ;
        RECT 5.295 0.085 5.545 0.885 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 4.560 1.105 4.730 1.275 ;
        RECT 4.920 1.105 5.090 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
      LAYER met1 ;
        RECT 3.465 1.305 4.105 1.320 ;
        RECT 3.465 1.075 5.150 1.305 ;
        RECT 3.465 1.060 4.105 1.075 ;
      LAYER via ;
        RECT 3.495 1.060 3.755 1.320 ;
        RECT 3.815 1.060 4.075 1.320 ;
      LAYER met2 ;
        RECT 3.445 1.005 4.125 1.375 ;
      LAYER via2 ;
        RECT 3.445 1.050 3.725 1.330 ;
        RECT 3.845 1.050 4.125 1.330 ;
      LAYER met3 ;
        RECT 3.395 1.025 4.175 1.355 ;
      LAYER via3 ;
        RECT 3.425 1.030 3.745 1.350 ;
        RECT 3.825 1.030 4.145 1.350 ;
      LAYER met4 ;
        RECT 1.370 0.680 4.150 1.860 ;
      LAYER via4 ;
        RECT 2.970 0.680 4.150 1.860 ;
      LAYER met5 ;
        RECT 1.250 0.560 4.270 1.945 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__probe_p_8

#--------EOF---------

MACRO sky130_fd_sc_hdll__probec_p_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__probec_p_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.832500 ;
    PORT
      LAYER li1 ;
        RECT 0.140 1.075 1.240 1.275 ;
    END
  END A
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 4.360 -0.155 6.675 0.560 ;
        RECT 4.560 -0.455 6.675 -0.155 ;
        RECT 4.360 -1.170 6.675 -0.455 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.635 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 4.360 3.175 6.675 3.890 ;
        RECT 4.560 2.875 6.675 3.175 ;
        RECT 4.360 2.160 6.675 2.875 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT -1.260 0.560 1.060 2.160 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.095 1.615 0.425 2.465 ;
        RECT 0.595 1.835 0.865 2.635 ;
        RECT 1.035 1.615 1.365 2.465 ;
        RECT 1.535 1.835 1.805 2.635 ;
        RECT 1.975 1.615 2.305 2.465 ;
        RECT 2.475 1.835 2.745 2.635 ;
        RECT 2.915 1.615 3.245 2.465 ;
        RECT 3.415 1.835 3.685 2.635 ;
        RECT 3.855 1.615 4.185 2.465 ;
        RECT 4.355 1.835 4.625 2.635 ;
        RECT 4.795 1.615 5.125 2.465 ;
        RECT 0.095 1.445 1.595 1.615 ;
        RECT 1.975 1.445 5.125 1.615 ;
        RECT 5.295 1.485 5.595 2.635 ;
        RECT 1.420 1.245 1.595 1.445 ;
        RECT 1.420 1.075 4.045 1.245 ;
        RECT 1.420 0.905 1.595 1.075 ;
        RECT 4.290 0.905 5.125 1.445 ;
        RECT 0.145 0.735 1.595 0.905 ;
        RECT 1.975 0.735 5.125 0.905 ;
        RECT 0.145 0.255 0.445 0.735 ;
        RECT 0.615 0.085 0.895 0.565 ;
        RECT 1.065 0.255 1.335 0.735 ;
        RECT 1.505 0.085 1.805 0.565 ;
        RECT 1.975 0.255 2.305 0.735 ;
        RECT 2.475 0.085 2.745 0.565 ;
        RECT 2.915 0.255 3.245 0.735 ;
        RECT 3.415 0.085 3.685 0.565 ;
        RECT 3.855 0.255 4.185 0.735 ;
        RECT 4.355 0.085 4.625 0.565 ;
        RECT 4.795 0.255 5.125 0.735 ;
        RECT 5.295 0.085 5.545 0.885 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 4.305 1.105 4.475 1.275 ;
        RECT 4.665 1.105 4.835 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
        RECT 2.020 1.260 2.660 1.320 ;
        RECT 4.245 1.260 4.895 1.305 ;
        RECT 2.020 1.120 4.895 1.260 ;
        RECT 2.020 1.060 2.660 1.120 ;
        RECT 4.245 1.075 4.895 1.120 ;
        RECT 0.000 -0.240 5.980 0.240 ;
      LAYER via ;
        RECT 5.230 2.590 5.490 2.850 ;
        RECT 5.550 2.590 5.810 2.850 ;
        RECT 2.050 1.060 2.310 1.320 ;
        RECT 2.370 1.060 2.630 1.320 ;
        RECT 5.230 -0.130 5.490 0.130 ;
        RECT 5.550 -0.130 5.810 0.130 ;
      LAYER met2 ;
        RECT 5.135 2.580 5.905 2.860 ;
        RECT 1.890 1.050 2.660 1.330 ;
        RECT 5.135 -0.140 5.905 0.140 ;
      LAYER via2 ;
        RECT 5.180 2.580 5.460 2.860 ;
        RECT 5.580 2.580 5.860 2.860 ;
        RECT 1.935 1.050 2.215 1.330 ;
        RECT 2.335 1.050 2.615 1.330 ;
        RECT 5.180 -0.140 5.460 0.140 ;
        RECT 5.580 -0.140 5.860 0.140 ;
      LAYER met3 ;
        RECT 5.130 2.555 5.910 2.885 ;
        RECT -0.715 1.030 0.065 1.350 ;
        RECT 1.885 1.025 2.665 1.355 ;
        RECT 5.130 -0.165 5.910 0.165 ;
      LAYER via3 ;
        RECT 5.160 2.560 5.480 2.880 ;
        RECT 5.560 2.560 5.880 2.880 ;
        RECT -0.685 1.030 -0.365 1.350 ;
        RECT -0.285 1.030 0.035 1.350 ;
        RECT 1.915 1.030 2.235 1.350 ;
        RECT 2.315 1.030 2.635 1.350 ;
        RECT 5.160 -0.160 5.480 0.160 ;
        RECT 5.560 -0.160 5.880 0.160 ;
      LAYER met4 ;
        RECT 4.930 2.435 6.110 3.615 ;
        RECT -1.140 0.770 0.040 1.950 ;
        RECT 1.460 0.770 2.640 1.950 ;
        RECT 4.930 -0.895 6.110 0.285 ;
      LAYER met5 ;
        RECT 1.160 -1.105 2.760 3.825 ;
        RECT 4.360 2.975 4.460 3.075 ;
        RECT 4.360 -0.355 4.460 -0.255 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__probec_p_8

#--------EOF---------

MACRO sky130_fd_sc_hdll__sdfbbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sdfbbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.640 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.435 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138600 ;
    PORT
      LAYER li1 ;
        RECT 4.155 1.325 4.475 2.375 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 12.515 1.095 13.090 1.325 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 1.490 1.025 1.765 1.685 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277200 ;
    PORT
      LAYER li1 ;
        RECT 1.935 1.015 2.255 1.695 ;
        RECT 1.935 0.765 2.605 1.015 ;
        RECT 1.935 0.760 2.255 0.765 ;
        RECT 1.975 0.345 2.255 0.760 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277200 ;
    PORT
      LAYER met1 ;
        RECT 6.525 0.920 6.815 0.965 ;
        RECT 10.655 0.920 10.945 0.965 ;
        RECT 6.525 0.780 10.945 0.920 ;
        RECT 6.525 0.735 6.815 0.780 ;
        RECT 10.655 0.735 10.945 0.780 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 15.640 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 13.010 1.005 15.600 1.015 ;
        RECT 6.750 0.785 9.225 1.005 ;
        RECT 11.025 0.785 15.600 1.005 ;
        RECT 0.005 0.105 15.600 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 15.830 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 15.640 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 15.260 1.605 15.545 2.465 ;
        RECT 15.310 0.825 15.545 1.605 ;
        RECT 15.260 0.255 15.545 0.825 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.595750 ;
    PORT
      LAYER li1 ;
        RECT 13.715 1.630 14.095 2.465 ;
        RECT 13.820 1.520 14.095 1.630 ;
        RECT 13.820 0.715 14.115 1.520 ;
        RECT 13.715 0.255 14.115 0.715 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 15.640 2.805 ;
        RECT 0.170 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.895 2.635 ;
        RECT 0.170 1.795 0.885 1.965 ;
        RECT 0.655 0.805 0.885 1.795 ;
        RECT 0.170 0.635 0.885 0.805 ;
        RECT 0.170 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.115 0.345 1.320 2.465 ;
        RECT 1.555 1.885 1.885 2.635 ;
        RECT 2.385 1.875 2.765 2.385 ;
        RECT 3.095 1.905 3.265 2.465 ;
        RECT 3.510 2.215 3.890 2.635 ;
        RECT 2.550 1.365 2.765 1.875 ;
        RECT 2.945 1.745 3.265 1.905 ;
        RECT 2.945 1.575 3.895 1.745 ;
        RECT 2.550 1.185 3.275 1.365 ;
        RECT 2.785 1.075 3.275 1.185 ;
        RECT 3.725 1.095 3.895 1.575 ;
        RECT 1.555 0.085 1.805 0.635 ;
        RECT 2.785 0.595 2.955 1.075 ;
        RECT 3.725 0.795 4.070 1.095 ;
        RECT 2.550 0.265 2.955 0.595 ;
        RECT 3.125 0.765 4.070 0.795 ;
        RECT 3.125 0.625 3.895 0.765 ;
        RECT 3.125 0.305 3.325 0.625 ;
        RECT 3.620 0.085 3.950 0.445 ;
        RECT 4.645 0.305 4.815 2.465 ;
        RECT 5.035 2.250 5.915 2.420 ;
        RECT 4.985 1.575 5.575 1.955 ;
        RECT 4.985 0.705 5.245 1.575 ;
        RECT 5.745 1.405 5.915 2.250 ;
        RECT 6.205 2.205 6.585 2.635 ;
        RECT 6.935 2.035 7.105 2.375 ;
        RECT 6.085 1.785 7.585 2.035 ;
        RECT 7.825 1.915 8.155 2.635 ;
        RECT 9.300 2.250 10.230 2.420 ;
        RECT 10.520 2.255 10.900 2.635 ;
        RECT 6.085 1.575 6.385 1.785 ;
        RECT 6.945 1.405 7.195 1.485 ;
        RECT 5.745 1.235 7.195 1.405 ;
        RECT 5.745 1.195 6.215 1.235 ;
        RECT 5.425 0.645 5.825 1.015 ;
        RECT 5.995 0.465 6.215 1.195 ;
        RECT 6.975 1.155 7.195 1.235 ;
        RECT 7.415 1.065 7.585 1.785 ;
        RECT 7.805 1.415 8.910 1.655 ;
        RECT 9.110 1.575 9.345 1.985 ;
        RECT 7.805 1.235 8.135 1.415 ;
        RECT 9.635 1.305 9.890 1.905 ;
        RECT 8.445 1.065 8.875 1.235 ;
        RECT 6.385 0.735 6.795 1.065 ;
        RECT 7.415 0.895 8.875 1.065 ;
        RECT 9.170 1.125 9.890 1.305 ;
        RECT 10.060 1.405 10.230 2.250 ;
        RECT 11.190 2.085 11.360 2.375 ;
        RECT 11.940 2.255 13.430 2.635 ;
        RECT 10.400 1.915 13.430 2.085 ;
        RECT 10.400 1.575 10.700 1.915 ;
        RECT 10.060 1.235 11.510 1.405 ;
        RECT 7.415 0.765 7.655 0.895 ;
        RECT 7.275 0.595 7.655 0.765 ;
        RECT 5.100 0.265 6.215 0.465 ;
        RECT 6.385 0.085 6.555 0.525 ;
        RECT 6.775 0.425 7.105 0.465 ;
        RECT 7.850 0.425 8.045 0.715 ;
        RECT 9.170 0.705 9.510 1.125 ;
        RECT 10.060 0.465 10.230 1.235 ;
        RECT 11.290 1.075 11.510 1.235 ;
        RECT 10.655 0.735 11.080 1.065 ;
        RECT 11.730 0.815 11.915 1.915 ;
        RECT 11.535 0.645 11.915 0.815 ;
        RECT 12.130 1.575 12.905 1.745 ;
        RECT 12.130 0.925 12.345 1.575 ;
        RECT 13.260 1.325 13.430 1.915 ;
        RECT 14.265 1.725 14.520 2.415 ;
        RECT 14.745 1.765 15.040 2.635 ;
        RECT 14.315 1.325 14.520 1.725 ;
        RECT 13.260 0.995 13.525 1.325 ;
        RECT 14.315 0.995 15.090 1.325 ;
        RECT 12.130 0.755 12.815 0.925 ;
        RECT 6.775 0.255 8.045 0.425 ;
        RECT 8.290 0.085 8.675 0.465 ;
        RECT 9.415 0.265 10.230 0.465 ;
        RECT 10.410 0.085 10.720 0.525 ;
        RECT 10.980 0.425 11.380 0.465 ;
        RECT 12.125 0.425 12.300 0.585 ;
        RECT 10.980 0.255 12.300 0.425 ;
        RECT 12.615 0.265 12.815 0.755 ;
        RECT 13.100 0.085 13.430 0.805 ;
        RECT 14.315 0.255 14.520 0.995 ;
        RECT 14.750 0.085 15.040 0.545 ;
        RECT 0.000 -0.085 15.640 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 14.405 2.635 14.575 2.805 ;
        RECT 14.865 2.635 15.035 2.805 ;
        RECT 15.325 2.635 15.495 2.805 ;
        RECT 0.655 1.785 0.825 1.955 ;
        RECT 1.150 0.765 1.320 0.935 ;
        RECT 3.105 1.105 3.275 1.275 ;
        RECT 4.645 1.105 4.815 1.275 ;
        RECT 5.145 1.785 5.315 1.955 ;
        RECT 5.655 0.765 5.825 0.935 ;
        RECT 9.175 1.785 9.345 1.955 ;
        RECT 8.715 1.445 8.885 1.615 ;
        RECT 6.585 0.765 6.755 0.935 ;
        RECT 9.175 1.105 9.345 1.275 ;
        RECT 10.715 0.765 10.885 0.935 ;
        RECT 12.165 1.445 12.335 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
        RECT 14.405 -0.085 14.575 0.085 ;
        RECT 14.865 -0.085 15.035 0.085 ;
        RECT 15.325 -0.085 15.495 0.085 ;
      LAYER met1 ;
        RECT 0.595 1.940 0.885 1.985 ;
        RECT 5.085 1.940 5.375 1.985 ;
        RECT 9.115 1.940 9.405 1.985 ;
        RECT 0.595 1.800 9.405 1.940 ;
        RECT 0.595 1.755 0.885 1.800 ;
        RECT 5.085 1.755 5.375 1.800 ;
        RECT 9.115 1.755 9.405 1.800 ;
        RECT 8.655 1.600 8.945 1.645 ;
        RECT 12.105 1.600 12.395 1.645 ;
        RECT 8.655 1.460 12.395 1.600 ;
        RECT 8.655 1.415 8.945 1.460 ;
        RECT 12.105 1.415 12.395 1.460 ;
        RECT 3.045 1.260 3.335 1.305 ;
        RECT 4.585 1.260 4.875 1.305 ;
        RECT 9.115 1.260 9.405 1.305 ;
        RECT 3.045 1.120 4.875 1.260 ;
        RECT 3.045 1.075 3.335 1.120 ;
        RECT 4.585 1.075 4.875 1.120 ;
        RECT 5.670 1.120 9.405 1.260 ;
        RECT 5.670 0.965 5.885 1.120 ;
        RECT 9.115 1.075 9.405 1.120 ;
        RECT 1.090 0.920 1.380 0.965 ;
        RECT 5.595 0.920 5.885 0.965 ;
        RECT 1.090 0.780 5.885 0.920 ;
        RECT 1.090 0.735 1.380 0.780 ;
        RECT 5.595 0.735 5.885 0.780 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfbbp_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__sdfrbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sdfrbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.260 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.140 0.975 0.490 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.160200 ;
    PORT
      LAYER li1 ;
        RECT 3.120 1.355 3.655 2.465 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277200 ;
    PORT
      LAYER met1 ;
        RECT 7.145 0.920 7.900 0.965 ;
        RECT 11.115 0.920 11.405 0.965 ;
        RECT 7.145 0.780 11.405 0.920 ;
        RECT 7.145 0.735 7.900 0.780 ;
        RECT 11.115 0.735 11.405 0.780 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.172800 ;
    PORT
      LAYER li1 ;
        RECT 4.610 0.710 4.955 1.700 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.467400 ;
    PORT
      LAYER li1 ;
        RECT 1.585 1.335 2.220 1.745 ;
        RECT 1.585 1.070 1.990 1.335 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 14.260 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.880 1.455 1.015 ;
        RECT 2.565 0.880 4.050 1.145 ;
        RECT 0.005 0.725 5.460 0.880 ;
        RECT 7.730 0.785 8.690 1.005 ;
        RECT 11.735 0.885 12.760 1.015 ;
        RECT 11.735 0.785 14.255 0.885 ;
        RECT 6.610 0.725 14.255 0.785 ;
        RECT 0.005 0.465 14.255 0.725 ;
        RECT 0.005 0.200 2.505 0.465 ;
        RECT 3.560 0.200 14.255 0.465 ;
        RECT 0.005 0.105 1.455 0.200 ;
        RECT 5.470 0.105 14.255 0.200 ;
        RECT 0.215 -0.010 0.235 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.425 14.450 2.910 ;
        RECT -0.190 1.305 2.120 1.425 ;
        RECT 4.455 1.305 14.450 1.425 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 14.260 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.513250 ;
    PORT
      LAYER li1 ;
        RECT 12.420 0.265 12.770 2.395 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.374700 ;
    PORT
      LAYER li1 ;
        RECT 13.885 1.475 14.165 2.465 ;
        RECT 13.935 0.870 14.165 1.475 ;
        RECT 13.885 0.255 14.165 0.870 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 14.260 2.805 ;
        RECT 0.090 1.965 0.345 2.465 ;
        RECT 0.530 2.135 0.910 2.635 ;
        RECT 0.090 1.795 0.915 1.965 ;
        RECT 0.710 1.325 0.915 1.795 ;
        RECT 1.135 1.730 1.365 2.465 ;
        RECT 2.110 2.085 2.380 2.400 ;
        RECT 2.600 2.255 2.930 2.635 ;
        RECT 3.870 2.105 4.040 2.465 ;
        RECT 4.855 2.275 5.205 2.635 ;
        RECT 5.480 2.185 5.850 2.435 ;
        RECT 5.480 2.105 5.650 2.185 ;
        RECT 6.095 2.135 6.460 2.465 ;
        RECT 2.110 1.915 2.730 2.085 ;
        RECT 0.710 0.995 1.025 1.325 ;
        RECT 0.710 0.805 0.885 0.995 ;
        RECT 0.095 0.635 0.885 0.805 ;
        RECT 1.195 0.675 1.365 1.730 ;
        RECT 2.475 1.185 2.730 1.915 ;
        RECT 3.870 1.935 5.650 2.105 ;
        RECT 2.475 1.165 3.445 1.185 ;
        RECT 2.265 0.995 3.445 1.165 ;
        RECT 3.870 1.075 4.045 1.935 ;
        RECT 2.265 0.900 2.435 0.995 ;
        RECT 0.095 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.115 0.345 1.365 0.675 ;
        RECT 1.695 0.730 2.435 0.900 ;
        RECT 1.695 0.395 1.865 0.730 ;
        RECT 2.035 0.085 2.415 0.560 ;
        RECT 2.655 0.085 3.035 0.825 ;
        RECT 3.275 0.425 3.445 0.995 ;
        RECT 3.665 0.675 4.045 1.075 ;
        RECT 4.265 0.425 4.435 1.685 ;
        RECT 5.140 0.895 5.310 1.935 ;
        RECT 5.820 1.575 6.120 1.955 ;
        RECT 5.480 1.065 5.650 1.395 ;
        RECT 5.900 1.035 6.120 1.575 ;
        RECT 6.290 1.385 6.460 2.135 ;
        RECT 6.680 2.105 6.850 2.375 ;
        RECT 7.135 2.355 7.465 2.635 ;
        RECT 7.770 2.105 7.940 2.375 ;
        RECT 8.150 2.175 8.570 2.635 ;
        RECT 6.680 1.935 7.940 2.105 ;
        RECT 8.815 2.005 8.985 2.465 ;
        RECT 9.195 2.125 10.215 2.465 ;
        RECT 10.415 2.195 10.665 2.635 ;
        RECT 8.230 1.835 8.985 2.005 ;
        RECT 8.230 1.765 8.540 1.835 ;
        RECT 6.960 1.595 8.540 1.765 ;
        RECT 9.185 1.665 9.845 1.955 ;
        RECT 6.290 1.215 8.150 1.385 ;
        RECT 5.140 0.715 5.720 0.895 ;
        RECT 3.275 0.255 4.435 0.425 ;
        RECT 5.005 0.085 5.350 0.540 ;
        RECT 5.550 0.505 5.720 0.715 ;
        RECT 5.900 0.705 6.650 1.035 ;
        RECT 5.550 0.335 5.890 0.505 ;
        RECT 6.840 0.475 7.010 1.215 ;
        RECT 7.230 0.765 7.810 1.045 ;
        RECT 7.980 1.005 8.150 1.215 ;
        RECT 8.370 0.835 8.540 1.595 ;
        RECT 6.110 0.305 7.010 0.475 ;
        RECT 7.690 0.085 8.020 0.545 ;
        RECT 8.230 0.445 8.540 0.835 ;
        RECT 8.710 1.660 9.845 1.665 ;
        RECT 10.040 1.745 10.215 2.125 ;
        RECT 10.910 2.085 11.080 2.375 ;
        RECT 11.255 2.255 11.635 2.635 ;
        RECT 10.910 1.915 11.730 2.085 ;
        RECT 8.710 1.495 9.445 1.660 ;
        RECT 10.040 1.575 11.370 1.745 ;
        RECT 8.710 0.705 8.970 1.495 ;
        RECT 10.040 1.485 10.285 1.575 ;
        RECT 9.235 0.920 9.405 1.325 ;
        RECT 9.670 1.315 10.285 1.485 ;
        RECT 11.560 1.325 11.730 1.915 ;
        RECT 11.905 1.495 12.190 2.635 ;
        RECT 12.940 1.705 13.110 2.465 ;
        RECT 13.285 1.875 13.695 2.635 ;
        RECT 12.940 1.535 13.605 1.705 ;
        RECT 13.435 1.325 13.605 1.535 ;
        RECT 9.670 0.535 9.890 1.315 ;
        RECT 10.150 0.865 10.370 1.145 ;
        RECT 10.600 1.065 11.370 1.275 ;
        RECT 10.150 0.695 10.730 0.865 ;
        RECT 8.230 0.275 8.610 0.445 ;
        RECT 8.780 0.255 9.890 0.535 ;
        RECT 10.110 0.085 10.330 0.525 ;
        RECT 10.560 0.465 10.730 0.695 ;
        RECT 11.065 0.635 11.370 1.065 ;
        RECT 11.560 0.995 12.205 1.325 ;
        RECT 13.435 0.995 13.765 1.325 ;
        RECT 11.560 0.465 11.735 0.995 ;
        RECT 13.435 0.805 13.605 0.995 ;
        RECT 10.560 0.295 11.735 0.465 ;
        RECT 11.905 0.085 12.190 0.710 ;
        RECT 12.940 0.635 13.605 0.805 ;
        RECT 12.940 0.255 13.110 0.635 ;
        RECT 13.285 0.085 13.695 0.465 ;
        RECT 0.000 -0.085 14.260 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 1.135 1.785 1.305 1.955 ;
        RECT 0.855 1.105 1.025 1.275 ;
        RECT 5.950 1.785 6.120 1.955 ;
        RECT 5.480 1.105 5.650 1.275 ;
        RECT 9.565 1.785 9.735 1.955 ;
        RECT 7.255 0.765 7.425 0.935 ;
        RECT 7.615 0.765 7.785 0.935 ;
        RECT 9.235 1.105 9.405 1.275 ;
        RECT 11.175 0.765 11.345 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
      LAYER met1 ;
        RECT 1.070 1.940 1.370 1.985 ;
        RECT 5.890 1.940 6.180 1.985 ;
        RECT 9.500 1.940 9.795 1.985 ;
        RECT 1.070 1.800 9.795 1.940 ;
        RECT 1.070 1.755 1.370 1.800 ;
        RECT 5.890 1.755 6.180 1.800 ;
        RECT 9.500 1.755 9.795 1.800 ;
        RECT 0.795 1.260 1.085 1.305 ;
        RECT 5.420 1.260 5.710 1.305 ;
        RECT 9.155 1.260 9.465 1.305 ;
        RECT 0.795 1.120 9.465 1.260 ;
        RECT 0.795 1.075 1.085 1.120 ;
        RECT 5.420 1.075 5.710 1.120 ;
        RECT 9.155 1.075 9.465 1.120 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfrbp_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__sdfrbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sdfrbp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.720 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.140 0.975 0.490 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.160200 ;
    PORT
      LAYER li1 ;
        RECT 3.120 1.355 3.655 2.465 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277200 ;
    PORT
      LAYER met1 ;
        RECT 7.145 0.920 7.900 0.965 ;
        RECT 11.115 0.920 11.405 0.965 ;
        RECT 7.145 0.780 11.405 0.920 ;
        RECT 7.145 0.735 7.900 0.780 ;
        RECT 11.115 0.735 11.405 0.780 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.172800 ;
    PORT
      LAYER li1 ;
        RECT 4.610 0.710 4.955 1.700 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.467400 ;
    PORT
      LAYER li1 ;
        RECT 1.585 1.335 2.220 1.745 ;
        RECT 1.585 1.070 1.990 1.335 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 14.720 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.880 1.455 1.015 ;
        RECT 2.565 0.880 4.050 1.145 ;
        RECT 0.005 0.725 5.460 0.880 ;
        RECT 7.730 0.785 8.690 1.005 ;
        RECT 12.265 0.785 14.715 1.015 ;
        RECT 6.610 0.725 14.715 0.785 ;
        RECT 0.005 0.465 14.715 0.725 ;
        RECT 0.005 0.200 2.505 0.465 ;
        RECT 3.560 0.200 14.715 0.465 ;
        RECT 0.005 0.105 1.455 0.200 ;
        RECT 5.470 0.105 14.715 0.200 ;
        RECT 0.215 -0.010 0.235 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.425 14.910 2.910 ;
        RECT -0.190 1.305 2.120 1.425 ;
        RECT 4.455 1.305 14.910 1.425 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 14.720 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.564000 ;
    PORT
      LAYER li1 ;
        RECT 12.860 0.265 13.260 1.695 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.494750 ;
    PORT
      LAYER li1 ;
        RECT 13.770 1.535 14.205 2.080 ;
        RECT 14.035 0.825 14.205 1.535 ;
        RECT 13.780 0.310 14.205 0.825 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 14.720 2.805 ;
        RECT 0.090 1.965 0.345 2.465 ;
        RECT 0.530 2.135 0.910 2.635 ;
        RECT 0.090 1.795 0.915 1.965 ;
        RECT 0.710 1.325 0.915 1.795 ;
        RECT 1.135 1.730 1.365 2.465 ;
        RECT 2.110 2.085 2.380 2.400 ;
        RECT 2.600 2.255 2.930 2.635 ;
        RECT 3.870 2.105 4.040 2.465 ;
        RECT 4.855 2.275 5.205 2.635 ;
        RECT 5.480 2.185 5.850 2.435 ;
        RECT 5.480 2.105 5.650 2.185 ;
        RECT 6.095 2.135 6.460 2.465 ;
        RECT 2.110 1.915 2.730 2.085 ;
        RECT 0.710 0.995 1.025 1.325 ;
        RECT 0.710 0.805 0.885 0.995 ;
        RECT 0.095 0.635 0.885 0.805 ;
        RECT 1.195 0.675 1.365 1.730 ;
        RECT 2.475 1.185 2.730 1.915 ;
        RECT 3.870 1.935 5.650 2.105 ;
        RECT 2.475 1.165 3.445 1.185 ;
        RECT 2.265 0.995 3.445 1.165 ;
        RECT 3.870 1.075 4.045 1.935 ;
        RECT 2.265 0.900 2.435 0.995 ;
        RECT 0.095 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.115 0.345 1.365 0.675 ;
        RECT 1.695 0.730 2.435 0.900 ;
        RECT 1.695 0.395 1.865 0.730 ;
        RECT 2.035 0.085 2.415 0.560 ;
        RECT 2.655 0.085 3.035 0.825 ;
        RECT 3.275 0.425 3.445 0.995 ;
        RECT 3.665 0.675 4.045 1.075 ;
        RECT 4.265 0.425 4.435 1.685 ;
        RECT 5.140 0.895 5.310 1.935 ;
        RECT 5.820 1.575 6.120 1.955 ;
        RECT 5.480 1.065 5.650 1.395 ;
        RECT 5.900 1.035 6.120 1.575 ;
        RECT 6.290 1.385 6.460 2.135 ;
        RECT 6.680 2.105 6.850 2.375 ;
        RECT 7.135 2.355 7.465 2.635 ;
        RECT 7.770 2.105 7.940 2.375 ;
        RECT 8.150 2.175 8.570 2.635 ;
        RECT 6.680 1.935 7.940 2.105 ;
        RECT 8.815 2.005 8.985 2.465 ;
        RECT 9.195 2.125 10.215 2.465 ;
        RECT 10.415 2.195 10.665 2.635 ;
        RECT 8.230 1.835 8.985 2.005 ;
        RECT 8.230 1.765 8.540 1.835 ;
        RECT 6.960 1.595 8.540 1.765 ;
        RECT 9.185 1.665 9.845 1.955 ;
        RECT 6.290 1.215 8.150 1.385 ;
        RECT 5.140 0.715 5.720 0.895 ;
        RECT 3.275 0.255 4.435 0.425 ;
        RECT 5.005 0.085 5.350 0.540 ;
        RECT 5.550 0.505 5.720 0.715 ;
        RECT 5.900 0.705 6.650 1.035 ;
        RECT 5.550 0.335 5.890 0.505 ;
        RECT 6.840 0.475 7.010 1.215 ;
        RECT 7.230 0.765 7.810 1.045 ;
        RECT 7.980 1.005 8.150 1.215 ;
        RECT 8.370 0.835 8.540 1.595 ;
        RECT 6.110 0.305 7.010 0.475 ;
        RECT 7.690 0.085 8.020 0.545 ;
        RECT 8.230 0.445 8.540 0.835 ;
        RECT 8.710 1.660 9.845 1.665 ;
        RECT 10.040 1.745 10.215 2.125 ;
        RECT 10.910 2.085 11.080 2.375 ;
        RECT 11.255 2.255 11.635 2.635 ;
        RECT 10.910 1.915 11.730 2.085 ;
        RECT 8.710 1.495 9.445 1.660 ;
        RECT 10.040 1.575 11.370 1.745 ;
        RECT 8.710 0.705 8.970 1.495 ;
        RECT 10.040 1.485 10.285 1.575 ;
        RECT 9.235 0.920 9.405 1.325 ;
        RECT 9.670 1.315 10.285 1.485 ;
        RECT 11.560 1.325 11.730 1.915 ;
        RECT 11.900 2.035 12.075 2.465 ;
        RECT 12.255 2.205 12.715 2.635 ;
        RECT 13.270 2.255 13.725 2.635 ;
        RECT 11.900 1.865 13.600 2.035 ;
        RECT 11.900 1.795 12.640 1.865 ;
        RECT 9.670 0.535 9.890 1.315 ;
        RECT 10.150 0.865 10.370 1.145 ;
        RECT 10.600 1.065 11.370 1.275 ;
        RECT 10.150 0.695 10.730 0.865 ;
        RECT 8.230 0.275 8.610 0.445 ;
        RECT 8.780 0.255 9.890 0.535 ;
        RECT 10.110 0.085 10.330 0.525 ;
        RECT 10.560 0.465 10.730 0.695 ;
        RECT 11.065 0.635 11.370 1.065 ;
        RECT 11.560 0.995 12.205 1.325 ;
        RECT 11.560 0.465 11.730 0.995 ;
        RECT 12.465 0.825 12.640 1.795 ;
        RECT 13.430 1.325 13.600 1.865 ;
        RECT 14.375 1.495 14.625 2.635 ;
        RECT 13.430 0.995 13.865 1.325 ;
        RECT 10.560 0.295 11.730 0.465 ;
        RECT 11.900 0.655 12.640 0.825 ;
        RECT 11.900 0.345 12.070 0.655 ;
        RECT 12.325 0.085 12.655 0.485 ;
        RECT 13.440 0.085 13.610 0.825 ;
        RECT 14.375 0.085 14.545 0.930 ;
        RECT 0.000 -0.085 14.720 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 14.405 2.635 14.575 2.805 ;
        RECT 1.135 1.785 1.305 1.955 ;
        RECT 0.855 1.105 1.025 1.275 ;
        RECT 5.950 1.785 6.120 1.955 ;
        RECT 5.480 1.105 5.650 1.275 ;
        RECT 9.565 1.785 9.735 1.955 ;
        RECT 7.255 0.765 7.425 0.935 ;
        RECT 7.615 0.765 7.785 0.935 ;
        RECT 9.235 1.105 9.405 1.275 ;
        RECT 11.175 0.765 11.345 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
        RECT 14.405 -0.085 14.575 0.085 ;
      LAYER met1 ;
        RECT 1.070 1.940 1.370 1.985 ;
        RECT 5.890 1.940 6.180 1.985 ;
        RECT 9.500 1.940 9.795 1.985 ;
        RECT 1.070 1.800 9.795 1.940 ;
        RECT 1.070 1.755 1.370 1.800 ;
        RECT 5.890 1.755 6.180 1.800 ;
        RECT 9.500 1.755 9.795 1.800 ;
        RECT 0.795 1.260 1.085 1.305 ;
        RECT 5.420 1.260 5.710 1.305 ;
        RECT 9.155 1.260 9.465 1.305 ;
        RECT 0.795 1.120 9.465 1.260 ;
        RECT 0.795 1.075 1.085 1.120 ;
        RECT 5.420 1.075 5.710 1.120 ;
        RECT 9.155 1.075 9.465 1.120 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfrbp_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__sdfrtn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sdfrtn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.880 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.140 0.975 0.490 1.625 ;
    END
  END CLK_N
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.160200 ;
    PORT
      LAYER li1 ;
        RECT 3.120 1.355 3.655 2.465 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277200 ;
    PORT
      LAYER met1 ;
        RECT 7.145 0.920 7.900 0.965 ;
        RECT 11.115 0.920 11.405 0.965 ;
        RECT 7.145 0.780 11.405 0.920 ;
        RECT 7.145 0.735 7.900 0.780 ;
        RECT 11.115 0.735 11.405 0.780 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.172800 ;
    PORT
      LAYER li1 ;
        RECT 4.610 0.710 4.955 1.700 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.467400 ;
    PORT
      LAYER li1 ;
        RECT 1.585 1.335 2.220 1.745 ;
        RECT 1.585 1.070 1.990 1.335 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 12.880 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.880 1.455 1.015 ;
        RECT 2.565 0.880 4.050 1.145 ;
        RECT 0.005 0.725 5.460 0.880 ;
        RECT 7.730 0.785 8.690 1.005 ;
        RECT 11.735 0.785 12.760 1.015 ;
        RECT 6.610 0.725 12.760 0.785 ;
        RECT 0.005 0.465 12.760 0.725 ;
        RECT 0.005 0.200 2.505 0.465 ;
        RECT 3.560 0.200 12.760 0.465 ;
        RECT 0.005 0.105 1.455 0.200 ;
        RECT 5.470 0.105 12.760 0.200 ;
        RECT 0.215 -0.010 0.235 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.425 13.070 2.910 ;
        RECT -0.190 1.305 2.120 1.425 ;
        RECT 4.455 1.305 13.070 1.425 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 12.880 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.513250 ;
    PORT
      LAYER li1 ;
        RECT 12.420 0.265 12.785 2.325 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 12.880 2.805 ;
        RECT 0.090 1.965 0.345 2.465 ;
        RECT 0.530 2.135 0.910 2.635 ;
        RECT 0.090 1.795 0.915 1.965 ;
        RECT 0.710 1.325 0.915 1.795 ;
        RECT 1.135 1.730 1.365 2.465 ;
        RECT 2.110 2.085 2.380 2.400 ;
        RECT 2.600 2.255 2.930 2.635 ;
        RECT 3.870 2.105 4.040 2.465 ;
        RECT 4.855 2.275 5.205 2.635 ;
        RECT 5.480 2.185 5.850 2.435 ;
        RECT 5.480 2.105 5.650 2.185 ;
        RECT 6.095 2.135 6.460 2.465 ;
        RECT 2.110 1.915 2.730 2.085 ;
        RECT 0.710 0.995 1.025 1.325 ;
        RECT 0.710 0.805 0.885 0.995 ;
        RECT 0.095 0.635 0.885 0.805 ;
        RECT 1.195 0.675 1.365 1.730 ;
        RECT 2.475 1.185 2.730 1.915 ;
        RECT 3.870 1.935 5.650 2.105 ;
        RECT 2.475 1.165 3.445 1.185 ;
        RECT 2.265 0.995 3.445 1.165 ;
        RECT 3.870 1.075 4.045 1.935 ;
        RECT 2.265 0.900 2.435 0.995 ;
        RECT 0.095 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.115 0.345 1.365 0.675 ;
        RECT 1.695 0.730 2.435 0.900 ;
        RECT 1.695 0.395 1.865 0.730 ;
        RECT 2.035 0.085 2.415 0.560 ;
        RECT 2.655 0.085 3.035 0.825 ;
        RECT 3.275 0.425 3.445 0.995 ;
        RECT 3.665 0.675 4.045 1.075 ;
        RECT 4.265 0.425 4.435 1.685 ;
        RECT 5.140 0.895 5.310 1.935 ;
        RECT 5.820 1.575 6.120 1.955 ;
        RECT 5.480 1.065 5.650 1.395 ;
        RECT 5.900 1.035 6.120 1.575 ;
        RECT 6.290 1.385 6.460 2.135 ;
        RECT 6.680 2.105 6.850 2.375 ;
        RECT 7.135 2.355 7.465 2.635 ;
        RECT 7.770 2.105 7.940 2.375 ;
        RECT 8.150 2.175 8.570 2.635 ;
        RECT 6.680 1.935 7.940 2.105 ;
        RECT 8.815 2.005 8.985 2.465 ;
        RECT 9.195 2.125 10.215 2.465 ;
        RECT 10.415 2.195 10.665 2.635 ;
        RECT 8.230 1.835 8.985 2.005 ;
        RECT 8.230 1.765 8.540 1.835 ;
        RECT 6.960 1.595 8.540 1.765 ;
        RECT 9.185 1.665 9.845 1.955 ;
        RECT 6.290 1.215 8.150 1.385 ;
        RECT 5.140 0.715 5.720 0.895 ;
        RECT 3.275 0.255 4.435 0.425 ;
        RECT 5.005 0.085 5.350 0.540 ;
        RECT 5.550 0.505 5.720 0.715 ;
        RECT 5.900 0.705 6.650 1.035 ;
        RECT 5.550 0.335 5.890 0.505 ;
        RECT 6.840 0.475 7.010 1.215 ;
        RECT 7.230 0.765 7.810 1.045 ;
        RECT 7.980 1.005 8.150 1.215 ;
        RECT 8.370 0.835 8.540 1.595 ;
        RECT 6.110 0.305 7.010 0.475 ;
        RECT 7.690 0.085 8.020 0.545 ;
        RECT 8.230 0.445 8.540 0.835 ;
        RECT 8.710 1.660 9.845 1.665 ;
        RECT 10.040 1.745 10.215 2.125 ;
        RECT 10.910 2.085 11.080 2.375 ;
        RECT 11.255 2.255 11.635 2.635 ;
        RECT 10.910 1.915 11.730 2.085 ;
        RECT 8.710 1.495 9.445 1.660 ;
        RECT 10.040 1.575 11.370 1.745 ;
        RECT 8.710 0.705 8.970 1.495 ;
        RECT 10.040 1.485 10.285 1.575 ;
        RECT 9.235 0.920 9.405 1.325 ;
        RECT 9.670 1.315 10.285 1.485 ;
        RECT 11.560 1.325 11.730 1.915 ;
        RECT 11.905 1.495 12.190 2.635 ;
        RECT 9.670 0.535 9.890 1.315 ;
        RECT 10.150 0.865 10.370 1.145 ;
        RECT 10.600 1.065 11.370 1.275 ;
        RECT 10.150 0.695 10.730 0.865 ;
        RECT 8.230 0.275 8.610 0.445 ;
        RECT 8.780 0.255 9.890 0.535 ;
        RECT 10.110 0.085 10.330 0.525 ;
        RECT 10.560 0.465 10.730 0.695 ;
        RECT 11.065 0.635 11.370 1.065 ;
        RECT 11.560 0.995 12.205 1.325 ;
        RECT 11.560 0.465 11.735 0.995 ;
        RECT 10.560 0.295 11.735 0.465 ;
        RECT 11.905 0.085 12.190 0.710 ;
        RECT 0.000 -0.085 12.880 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 0.725 1.785 0.895 1.955 ;
        RECT 1.195 1.105 1.365 1.275 ;
        RECT 5.950 1.785 6.120 1.955 ;
        RECT 5.480 1.105 5.650 1.275 ;
        RECT 9.565 1.785 9.735 1.955 ;
        RECT 7.255 0.765 7.425 0.935 ;
        RECT 7.615 0.765 7.785 0.935 ;
        RECT 9.235 1.105 9.405 1.275 ;
        RECT 11.175 0.765 11.345 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
      LAYER met1 ;
        RECT 0.660 1.940 0.960 1.985 ;
        RECT 5.890 1.940 6.180 1.985 ;
        RECT 9.500 1.940 9.795 1.985 ;
        RECT 0.660 1.800 9.795 1.940 ;
        RECT 0.660 1.755 0.960 1.800 ;
        RECT 5.890 1.755 6.180 1.800 ;
        RECT 9.500 1.755 9.795 1.800 ;
        RECT 1.135 1.260 1.425 1.305 ;
        RECT 5.420 1.260 5.710 1.305 ;
        RECT 9.155 1.260 9.465 1.305 ;
        RECT 1.135 1.120 9.465 1.260 ;
        RECT 1.135 1.075 1.425 1.120 ;
        RECT 5.420 1.075 5.710 1.120 ;
        RECT 9.155 1.075 9.465 1.120 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfrtn_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__sdfrtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sdfrtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.880 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.140 0.975 0.490 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.160200 ;
    PORT
      LAYER li1 ;
        RECT 3.120 1.355 3.655 2.465 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277200 ;
    PORT
      LAYER met1 ;
        RECT 7.145 0.920 7.900 0.965 ;
        RECT 11.115 0.920 11.405 0.965 ;
        RECT 7.145 0.780 11.405 0.920 ;
        RECT 7.145 0.735 7.900 0.780 ;
        RECT 11.115 0.735 11.405 0.780 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.172800 ;
    PORT
      LAYER li1 ;
        RECT 4.610 0.710 4.955 1.700 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.467400 ;
    PORT
      LAYER li1 ;
        RECT 1.585 1.335 2.220 1.745 ;
        RECT 1.585 1.070 1.990 1.335 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 12.880 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.880 1.455 1.015 ;
        RECT 2.565 0.880 4.050 1.145 ;
        RECT 0.005 0.725 5.460 0.880 ;
        RECT 7.730 0.785 8.690 1.005 ;
        RECT 11.735 0.785 12.760 1.015 ;
        RECT 6.610 0.725 12.760 0.785 ;
        RECT 0.005 0.465 12.760 0.725 ;
        RECT 0.005 0.200 2.505 0.465 ;
        RECT 3.560 0.200 12.760 0.465 ;
        RECT 0.005 0.105 1.455 0.200 ;
        RECT 5.470 0.105 12.760 0.200 ;
        RECT 0.215 -0.010 0.235 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.425 13.070 2.910 ;
        RECT -0.190 1.305 2.120 1.425 ;
        RECT 4.455 1.305 13.070 1.425 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 12.880 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.513250 ;
    PORT
      LAYER li1 ;
        RECT 12.420 0.265 12.785 2.325 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 12.880 2.805 ;
        RECT 0.090 1.965 0.345 2.465 ;
        RECT 0.530 2.135 0.910 2.635 ;
        RECT 0.090 1.795 0.915 1.965 ;
        RECT 0.710 1.325 0.915 1.795 ;
        RECT 1.135 1.730 1.365 2.465 ;
        RECT 2.110 2.085 2.380 2.400 ;
        RECT 2.600 2.255 2.930 2.635 ;
        RECT 3.870 2.105 4.040 2.465 ;
        RECT 4.855 2.275 5.205 2.635 ;
        RECT 5.480 2.185 5.850 2.435 ;
        RECT 5.480 2.105 5.650 2.185 ;
        RECT 6.095 2.135 6.460 2.465 ;
        RECT 2.110 1.915 2.730 2.085 ;
        RECT 0.710 0.995 1.025 1.325 ;
        RECT 0.710 0.805 0.885 0.995 ;
        RECT 0.095 0.635 0.885 0.805 ;
        RECT 1.195 0.675 1.365 1.730 ;
        RECT 2.475 1.185 2.730 1.915 ;
        RECT 3.870 1.935 5.650 2.105 ;
        RECT 2.475 1.165 3.445 1.185 ;
        RECT 2.265 0.995 3.445 1.165 ;
        RECT 3.870 1.075 4.045 1.935 ;
        RECT 2.265 0.900 2.435 0.995 ;
        RECT 0.095 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.115 0.345 1.365 0.675 ;
        RECT 1.695 0.730 2.435 0.900 ;
        RECT 1.695 0.395 1.865 0.730 ;
        RECT 2.035 0.085 2.415 0.560 ;
        RECT 2.655 0.085 3.035 0.825 ;
        RECT 3.275 0.425 3.445 0.995 ;
        RECT 3.665 0.675 4.045 1.075 ;
        RECT 4.265 0.425 4.435 1.685 ;
        RECT 5.140 0.895 5.310 1.935 ;
        RECT 5.820 1.575 6.120 1.955 ;
        RECT 5.480 1.065 5.650 1.395 ;
        RECT 5.900 1.035 6.120 1.575 ;
        RECT 6.290 1.385 6.460 2.135 ;
        RECT 6.680 2.105 6.850 2.375 ;
        RECT 7.135 2.355 7.465 2.635 ;
        RECT 7.770 2.105 7.940 2.375 ;
        RECT 8.150 2.175 8.570 2.635 ;
        RECT 6.680 1.935 7.940 2.105 ;
        RECT 8.815 2.005 8.985 2.465 ;
        RECT 9.195 2.125 10.215 2.465 ;
        RECT 10.415 2.195 10.665 2.635 ;
        RECT 8.230 1.835 8.985 2.005 ;
        RECT 8.230 1.765 8.540 1.835 ;
        RECT 6.960 1.595 8.540 1.765 ;
        RECT 9.185 1.665 9.845 1.955 ;
        RECT 6.290 1.215 8.150 1.385 ;
        RECT 5.140 0.715 5.720 0.895 ;
        RECT 3.275 0.255 4.435 0.425 ;
        RECT 5.005 0.085 5.350 0.540 ;
        RECT 5.550 0.505 5.720 0.715 ;
        RECT 5.900 0.705 6.650 1.035 ;
        RECT 5.550 0.335 5.890 0.505 ;
        RECT 6.840 0.475 7.010 1.215 ;
        RECT 7.230 0.765 7.810 1.045 ;
        RECT 7.980 1.005 8.150 1.215 ;
        RECT 8.370 0.835 8.540 1.595 ;
        RECT 6.110 0.305 7.010 0.475 ;
        RECT 7.690 0.085 8.020 0.545 ;
        RECT 8.230 0.445 8.540 0.835 ;
        RECT 8.710 1.660 9.845 1.665 ;
        RECT 10.040 1.745 10.215 2.125 ;
        RECT 10.910 2.085 11.080 2.375 ;
        RECT 11.255 2.255 11.635 2.635 ;
        RECT 10.910 1.915 11.730 2.085 ;
        RECT 8.710 1.495 9.445 1.660 ;
        RECT 10.040 1.575 11.370 1.745 ;
        RECT 8.710 0.705 8.970 1.495 ;
        RECT 10.040 1.485 10.285 1.575 ;
        RECT 9.235 0.920 9.405 1.325 ;
        RECT 9.670 1.315 10.285 1.485 ;
        RECT 11.560 1.325 11.730 1.915 ;
        RECT 11.905 1.495 12.190 2.635 ;
        RECT 9.670 0.535 9.890 1.315 ;
        RECT 10.150 0.865 10.370 1.145 ;
        RECT 10.600 1.065 11.370 1.275 ;
        RECT 10.150 0.695 10.730 0.865 ;
        RECT 8.230 0.275 8.610 0.445 ;
        RECT 8.780 0.255 9.890 0.535 ;
        RECT 10.110 0.085 10.330 0.525 ;
        RECT 10.560 0.465 10.730 0.695 ;
        RECT 11.065 0.635 11.370 1.065 ;
        RECT 11.560 0.995 12.205 1.325 ;
        RECT 11.560 0.465 11.735 0.995 ;
        RECT 10.560 0.295 11.735 0.465 ;
        RECT 11.905 0.085 12.190 0.710 ;
        RECT 0.000 -0.085 12.880 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 1.135 1.785 1.305 1.955 ;
        RECT 0.855 1.105 1.025 1.275 ;
        RECT 5.950 1.785 6.120 1.955 ;
        RECT 5.480 1.105 5.650 1.275 ;
        RECT 9.565 1.785 9.735 1.955 ;
        RECT 7.255 0.765 7.425 0.935 ;
        RECT 7.615 0.765 7.785 0.935 ;
        RECT 9.235 1.105 9.405 1.275 ;
        RECT 11.175 0.765 11.345 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
      LAYER met1 ;
        RECT 1.070 1.940 1.370 1.985 ;
        RECT 5.890 1.940 6.180 1.985 ;
        RECT 9.500 1.940 9.795 1.985 ;
        RECT 1.070 1.800 9.795 1.940 ;
        RECT 1.070 1.755 1.370 1.800 ;
        RECT 5.890 1.755 6.180 1.800 ;
        RECT 9.500 1.755 9.795 1.800 ;
        RECT 0.795 1.260 1.085 1.305 ;
        RECT 5.420 1.260 5.710 1.305 ;
        RECT 9.155 1.260 9.465 1.305 ;
        RECT 0.795 1.120 9.465 1.260 ;
        RECT 0.795 1.075 1.085 1.120 ;
        RECT 5.420 1.075 5.710 1.120 ;
        RECT 9.155 1.075 9.465 1.120 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfrtp_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__sdfrtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sdfrtp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.340 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.140 0.975 0.490 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.160200 ;
    PORT
      LAYER li1 ;
        RECT 3.120 1.355 3.655 2.465 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277200 ;
    PORT
      LAYER met1 ;
        RECT 7.145 0.920 7.900 0.965 ;
        RECT 11.080 0.920 11.370 0.965 ;
        RECT 7.145 0.780 11.370 0.920 ;
        RECT 7.145 0.735 7.900 0.780 ;
        RECT 11.080 0.735 11.370 0.780 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.172800 ;
    PORT
      LAYER li1 ;
        RECT 4.610 0.710 4.955 1.700 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.467400 ;
    PORT
      LAYER li1 ;
        RECT 1.585 1.335 2.220 1.745 ;
        RECT 1.585 1.070 1.990 1.335 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 13.340 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.880 1.455 1.015 ;
        RECT 2.565 0.880 4.050 1.145 ;
        RECT 0.005 0.725 5.460 0.880 ;
        RECT 7.730 0.785 8.690 1.005 ;
        RECT 11.735 0.785 13.335 1.015 ;
        RECT 6.610 0.725 13.335 0.785 ;
        RECT 0.005 0.465 13.335 0.725 ;
        RECT 0.005 0.200 2.505 0.465 ;
        RECT 3.560 0.200 13.335 0.465 ;
        RECT 0.005 0.105 1.455 0.200 ;
        RECT 5.470 0.105 13.335 0.200 ;
        RECT 0.215 -0.010 0.235 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.425 13.530 2.910 ;
        RECT -0.190 1.305 2.120 1.425 ;
        RECT 4.455 1.305 13.530 1.425 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 13.340 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.498000 ;
    PORT
      LAYER li1 ;
        RECT 12.500 0.265 12.785 2.325 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 13.340 2.805 ;
        RECT 0.090 1.965 0.345 2.465 ;
        RECT 0.530 2.135 0.910 2.635 ;
        RECT 0.090 1.795 0.915 1.965 ;
        RECT 0.710 1.325 0.915 1.795 ;
        RECT 1.135 1.730 1.365 2.465 ;
        RECT 2.110 2.085 2.380 2.400 ;
        RECT 2.600 2.255 2.930 2.635 ;
        RECT 3.870 2.105 4.040 2.465 ;
        RECT 4.855 2.275 5.205 2.635 ;
        RECT 5.480 2.185 5.850 2.435 ;
        RECT 5.480 2.105 5.650 2.185 ;
        RECT 6.095 2.135 6.460 2.465 ;
        RECT 2.110 1.915 2.730 2.085 ;
        RECT 0.710 0.995 1.025 1.325 ;
        RECT 0.710 0.805 0.885 0.995 ;
        RECT 0.095 0.635 0.885 0.805 ;
        RECT 1.195 0.675 1.365 1.730 ;
        RECT 2.475 1.185 2.730 1.915 ;
        RECT 3.870 1.935 5.650 2.105 ;
        RECT 2.475 1.165 3.445 1.185 ;
        RECT 2.265 0.995 3.445 1.165 ;
        RECT 3.870 1.075 4.045 1.935 ;
        RECT 2.265 0.900 2.435 0.995 ;
        RECT 0.095 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.115 0.345 1.365 0.675 ;
        RECT 1.695 0.730 2.435 0.900 ;
        RECT 1.695 0.395 1.865 0.730 ;
        RECT 2.035 0.085 2.415 0.560 ;
        RECT 2.655 0.085 3.035 0.825 ;
        RECT 3.275 0.425 3.445 0.995 ;
        RECT 3.665 0.675 4.045 1.075 ;
        RECT 4.265 0.425 4.435 1.685 ;
        RECT 5.140 0.895 5.310 1.935 ;
        RECT 5.820 1.575 6.120 1.955 ;
        RECT 5.480 1.065 5.650 1.395 ;
        RECT 5.900 1.035 6.120 1.575 ;
        RECT 6.290 1.385 6.460 2.135 ;
        RECT 6.680 2.105 6.850 2.375 ;
        RECT 7.135 2.355 7.465 2.635 ;
        RECT 7.770 2.105 7.940 2.375 ;
        RECT 8.150 2.175 8.570 2.635 ;
        RECT 6.680 1.935 7.940 2.105 ;
        RECT 8.815 2.005 8.985 2.465 ;
        RECT 9.195 2.125 10.215 2.465 ;
        RECT 10.415 2.195 10.665 2.635 ;
        RECT 8.230 1.835 8.985 2.005 ;
        RECT 8.230 1.765 8.540 1.835 ;
        RECT 6.960 1.595 8.540 1.765 ;
        RECT 9.185 1.665 9.845 1.955 ;
        RECT 6.290 1.215 8.150 1.385 ;
        RECT 5.140 0.715 5.720 0.895 ;
        RECT 3.275 0.255 4.435 0.425 ;
        RECT 5.005 0.085 5.350 0.540 ;
        RECT 5.550 0.505 5.720 0.715 ;
        RECT 5.900 0.705 6.650 1.035 ;
        RECT 5.550 0.335 5.890 0.505 ;
        RECT 6.840 0.475 7.010 1.215 ;
        RECT 7.230 0.765 7.810 1.045 ;
        RECT 7.980 1.005 8.150 1.215 ;
        RECT 8.370 0.835 8.540 1.595 ;
        RECT 6.110 0.305 7.010 0.475 ;
        RECT 7.690 0.085 8.020 0.545 ;
        RECT 8.230 0.445 8.540 0.835 ;
        RECT 8.710 1.660 9.845 1.665 ;
        RECT 10.040 1.745 10.215 2.125 ;
        RECT 10.910 2.085 11.080 2.375 ;
        RECT 11.255 2.255 11.635 2.635 ;
        RECT 10.910 1.915 11.730 2.085 ;
        RECT 8.710 1.495 9.445 1.660 ;
        RECT 10.040 1.575 11.370 1.745 ;
        RECT 8.710 0.705 8.970 1.495 ;
        RECT 10.040 1.485 10.285 1.575 ;
        RECT 9.235 0.920 9.405 1.325 ;
        RECT 9.670 1.315 10.285 1.485 ;
        RECT 11.560 1.325 11.730 1.915 ;
        RECT 11.905 1.495 12.330 2.635 ;
        RECT 12.995 1.495 13.245 2.635 ;
        RECT 9.670 0.535 9.890 1.315 ;
        RECT 10.150 0.865 10.370 1.145 ;
        RECT 10.600 1.065 11.370 1.275 ;
        RECT 10.150 0.695 10.730 0.865 ;
        RECT 8.230 0.275 8.610 0.445 ;
        RECT 8.780 0.255 9.890 0.535 ;
        RECT 10.110 0.085 10.330 0.525 ;
        RECT 10.560 0.465 10.730 0.695 ;
        RECT 11.065 0.635 11.370 1.065 ;
        RECT 11.560 0.995 12.235 1.325 ;
        RECT 11.560 0.465 11.735 0.995 ;
        RECT 10.560 0.295 11.735 0.465 ;
        RECT 11.905 0.085 12.325 0.670 ;
        RECT 12.995 0.085 13.165 0.545 ;
        RECT 0.000 -0.085 13.340 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 1.135 1.785 1.305 1.955 ;
        RECT 0.855 1.105 1.025 1.275 ;
        RECT 5.950 1.785 6.120 1.955 ;
        RECT 5.480 1.105 5.650 1.275 ;
        RECT 9.565 1.785 9.735 1.955 ;
        RECT 7.255 0.765 7.425 0.935 ;
        RECT 7.615 0.765 7.785 0.935 ;
        RECT 9.235 1.105 9.405 1.275 ;
        RECT 11.140 0.765 11.310 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
      LAYER met1 ;
        RECT 1.070 1.940 1.370 1.985 ;
        RECT 5.890 1.940 6.180 1.985 ;
        RECT 9.500 1.940 9.795 1.985 ;
        RECT 1.070 1.800 9.795 1.940 ;
        RECT 1.070 1.755 1.370 1.800 ;
        RECT 5.890 1.755 6.180 1.800 ;
        RECT 9.500 1.755 9.795 1.800 ;
        RECT 0.795 1.260 1.085 1.305 ;
        RECT 5.420 1.260 5.710 1.305 ;
        RECT 9.155 1.260 9.465 1.305 ;
        RECT 0.795 1.120 9.465 1.260 ;
        RECT 0.795 1.075 1.085 1.120 ;
        RECT 5.420 1.075 5.710 1.120 ;
        RECT 9.155 1.075 9.465 1.120 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfrtp_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__sdfrtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sdfrtp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.260 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.140 0.975 0.490 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.160200 ;
    PORT
      LAYER li1 ;
        RECT 3.120 1.355 3.655 2.465 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277200 ;
    PORT
      LAYER met1 ;
        RECT 10.775 0.965 11.065 1.310 ;
        RECT 7.145 0.920 7.900 0.965 ;
        RECT 10.775 0.920 11.405 0.965 ;
        RECT 7.145 0.780 11.405 0.920 ;
        RECT 7.145 0.735 7.900 0.780 ;
        RECT 11.115 0.735 11.405 0.780 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.172800 ;
    PORT
      LAYER li1 ;
        RECT 4.610 0.710 4.955 1.700 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.467400 ;
    PORT
      LAYER li1 ;
        RECT 1.585 1.335 2.220 1.745 ;
        RECT 1.585 1.070 1.990 1.335 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 14.260 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.880 1.455 1.015 ;
        RECT 2.565 0.880 4.050 1.145 ;
        RECT 0.005 0.725 5.460 0.880 ;
        RECT 7.730 0.785 8.690 1.005 ;
        RECT 11.735 0.785 14.255 1.015 ;
        RECT 6.610 0.725 14.255 0.785 ;
        RECT 0.005 0.465 14.255 0.725 ;
        RECT 0.005 0.200 2.505 0.465 ;
        RECT 3.560 0.200 14.255 0.465 ;
        RECT 0.005 0.105 1.455 0.200 ;
        RECT 5.470 0.105 14.255 0.200 ;
        RECT 0.215 -0.010 0.235 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.425 14.450 2.910 ;
        RECT -0.190 1.305 2.120 1.425 ;
        RECT 4.455 1.305 14.450 1.425 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 14.260 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.171500 ;
    PORT
      LAYER li1 ;
        RECT 12.425 1.325 12.755 2.325 ;
        RECT 13.445 1.325 13.695 2.325 ;
        RECT 12.425 0.995 13.695 1.325 ;
        RECT 12.425 0.265 12.755 0.995 ;
        RECT 13.445 0.265 13.695 0.995 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 14.260 2.805 ;
        RECT 0.090 1.965 0.345 2.465 ;
        RECT 0.530 2.135 0.910 2.635 ;
        RECT 0.090 1.795 0.915 1.965 ;
        RECT 0.710 1.325 0.915 1.795 ;
        RECT 1.135 1.730 1.365 2.465 ;
        RECT 2.110 2.085 2.380 2.400 ;
        RECT 2.600 2.255 2.930 2.635 ;
        RECT 3.870 2.105 4.040 2.465 ;
        RECT 4.855 2.275 5.205 2.635 ;
        RECT 5.480 2.185 5.850 2.435 ;
        RECT 5.480 2.105 5.650 2.185 ;
        RECT 6.095 2.135 6.460 2.465 ;
        RECT 2.110 1.915 2.730 2.085 ;
        RECT 0.710 0.995 1.025 1.325 ;
        RECT 0.710 0.805 0.885 0.995 ;
        RECT 0.095 0.635 0.885 0.805 ;
        RECT 1.195 0.675 1.365 1.730 ;
        RECT 2.475 1.185 2.730 1.915 ;
        RECT 3.870 1.935 5.650 2.105 ;
        RECT 2.475 1.165 3.445 1.185 ;
        RECT 2.265 0.995 3.445 1.165 ;
        RECT 3.870 1.075 4.045 1.935 ;
        RECT 2.265 0.900 2.435 0.995 ;
        RECT 0.095 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.115 0.345 1.365 0.675 ;
        RECT 1.695 0.730 2.435 0.900 ;
        RECT 1.695 0.395 1.865 0.730 ;
        RECT 2.035 0.085 2.415 0.560 ;
        RECT 2.655 0.085 3.035 0.825 ;
        RECT 3.275 0.425 3.445 0.995 ;
        RECT 3.665 0.675 4.045 1.075 ;
        RECT 4.265 0.425 4.435 1.685 ;
        RECT 5.140 0.895 5.310 1.935 ;
        RECT 5.820 1.575 6.120 1.955 ;
        RECT 5.480 1.065 5.650 1.395 ;
        RECT 5.900 1.035 6.120 1.575 ;
        RECT 6.290 1.385 6.460 2.135 ;
        RECT 6.680 2.105 6.850 2.375 ;
        RECT 7.135 2.355 7.465 2.635 ;
        RECT 7.770 2.105 7.940 2.375 ;
        RECT 8.150 2.175 8.570 2.635 ;
        RECT 6.680 1.935 7.940 2.105 ;
        RECT 8.815 2.005 8.985 2.465 ;
        RECT 9.195 2.125 10.215 2.465 ;
        RECT 10.415 2.195 10.665 2.635 ;
        RECT 8.230 1.835 8.985 2.005 ;
        RECT 8.230 1.765 8.540 1.835 ;
        RECT 6.960 1.595 8.540 1.765 ;
        RECT 9.185 1.665 9.845 1.955 ;
        RECT 6.290 1.215 8.150 1.385 ;
        RECT 5.140 0.715 5.720 0.895 ;
        RECT 3.275 0.255 4.435 0.425 ;
        RECT 5.005 0.085 5.350 0.540 ;
        RECT 5.550 0.505 5.720 0.715 ;
        RECT 5.900 0.705 6.650 1.035 ;
        RECT 5.550 0.335 5.890 0.505 ;
        RECT 6.840 0.475 7.010 1.215 ;
        RECT 7.230 0.765 7.810 1.045 ;
        RECT 7.980 1.005 8.150 1.215 ;
        RECT 8.370 0.835 8.540 1.595 ;
        RECT 6.110 0.305 7.010 0.475 ;
        RECT 7.690 0.085 8.020 0.545 ;
        RECT 8.230 0.445 8.540 0.835 ;
        RECT 8.710 1.660 9.845 1.665 ;
        RECT 10.040 1.745 10.215 2.125 ;
        RECT 10.910 2.085 11.080 2.375 ;
        RECT 11.255 2.255 11.635 2.635 ;
        RECT 10.910 1.915 11.730 2.085 ;
        RECT 8.710 1.495 9.445 1.660 ;
        RECT 10.040 1.575 11.370 1.745 ;
        RECT 8.710 0.705 8.970 1.495 ;
        RECT 10.040 1.485 10.285 1.575 ;
        RECT 9.235 0.920 9.405 1.325 ;
        RECT 9.670 1.315 10.285 1.485 ;
        RECT 11.560 1.325 11.730 1.915 ;
        RECT 11.905 1.495 12.155 2.635 ;
        RECT 12.975 1.495 13.225 2.635 ;
        RECT 13.915 1.495 14.165 2.635 ;
        RECT 9.670 0.535 9.890 1.315 ;
        RECT 10.150 0.865 10.370 1.145 ;
        RECT 10.600 1.065 11.370 1.275 ;
        RECT 10.150 0.695 10.730 0.865 ;
        RECT 8.230 0.275 8.610 0.445 ;
        RECT 8.780 0.255 9.890 0.535 ;
        RECT 10.110 0.085 10.330 0.525 ;
        RECT 10.560 0.465 10.730 0.695 ;
        RECT 11.065 0.635 11.370 1.065 ;
        RECT 11.560 0.995 12.205 1.325 ;
        RECT 11.560 0.465 11.735 0.995 ;
        RECT 10.560 0.295 11.735 0.465 ;
        RECT 11.905 0.085 12.075 0.545 ;
        RECT 12.975 0.085 13.145 0.545 ;
        RECT 13.915 0.085 14.085 0.545 ;
        RECT 0.000 -0.085 14.260 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 1.135 1.785 1.305 1.955 ;
        RECT 0.855 1.105 1.025 1.275 ;
        RECT 5.950 1.785 6.120 1.955 ;
        RECT 5.480 1.105 5.650 1.275 ;
        RECT 9.565 1.785 9.735 1.955 ;
        RECT 7.255 0.765 7.425 0.935 ;
        RECT 7.615 0.765 7.785 0.935 ;
        RECT 9.235 1.105 9.405 1.275 ;
        RECT 10.835 1.085 11.005 1.255 ;
        RECT 11.175 0.765 11.345 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
      LAYER met1 ;
        RECT 1.070 1.940 1.370 1.985 ;
        RECT 5.890 1.940 6.180 1.985 ;
        RECT 9.500 1.940 9.795 1.985 ;
        RECT 1.070 1.800 9.795 1.940 ;
        RECT 1.070 1.755 1.370 1.800 ;
        RECT 5.890 1.755 6.180 1.800 ;
        RECT 9.500 1.755 9.795 1.800 ;
        RECT 0.795 1.260 1.085 1.305 ;
        RECT 5.420 1.260 5.710 1.305 ;
        RECT 9.155 1.260 9.465 1.305 ;
        RECT 0.795 1.120 9.465 1.260 ;
        RECT 0.795 1.075 1.085 1.120 ;
        RECT 5.420 1.075 5.710 1.120 ;
        RECT 9.155 1.075 9.465 1.120 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfrtp_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__sdfsbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sdfsbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.720 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 2.855 1.720 3.335 1.970 ;
        RECT 3.155 1.590 3.335 1.720 ;
        RECT 3.155 1.055 3.815 1.590 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 1.030 0.765 1.425 1.675 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.365 1.675 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.356400 ;
    PORT
      LAYER met1 ;
        RECT 0.570 1.260 0.860 1.305 ;
        RECT 2.585 1.260 2.875 1.305 ;
        RECT 0.570 1.120 2.875 1.260 ;
        RECT 0.570 1.075 0.860 1.120 ;
        RECT 2.585 1.075 2.875 1.120 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277200 ;
    PORT
      LAYER met1 ;
        RECT 7.385 1.600 7.725 1.645 ;
        RECT 9.675 1.600 9.965 1.645 ;
        RECT 7.385 1.460 9.965 1.600 ;
        RECT 7.385 1.415 7.725 1.460 ;
        RECT 9.675 1.415 9.965 1.460 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 14.720 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 7.690 0.785 9.595 1.005 ;
        RECT 12.040 0.785 14.535 1.015 ;
        RECT 0.005 0.105 14.535 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 14.910 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 14.720 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 14.065 1.495 14.625 2.450 ;
        RECT 14.270 0.825 14.625 1.495 ;
        RECT 14.065 0.275 14.625 0.825 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.471500 ;
    PORT
      LAYER li1 ;
        RECT 12.550 0.255 12.930 2.465 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 14.720 2.805 ;
        RECT 0.085 2.025 0.345 2.465 ;
        RECT 0.515 2.195 0.815 2.635 ;
        RECT 1.035 2.255 2.245 2.465 ;
        RECT 1.035 2.025 1.205 2.255 ;
        RECT 2.470 2.085 2.685 2.465 ;
        RECT 2.940 2.140 3.280 2.635 ;
        RECT 0.085 1.845 1.205 2.025 ;
        RECT 1.395 1.870 1.845 2.075 ;
        RECT 0.550 0.765 0.860 1.675 ;
        RECT 0.085 0.085 0.430 0.595 ;
        RECT 1.655 0.560 1.845 1.870 ;
        RECT 2.065 1.770 2.685 2.085 ;
        RECT 3.505 1.955 3.675 2.325 ;
        RECT 3.845 2.275 4.225 2.635 ;
        RECT 4.445 2.135 4.790 2.465 ;
        RECT 3.505 1.775 4.295 1.955 ;
        RECT 2.065 0.905 2.400 1.770 ;
        RECT 2.570 1.075 2.950 1.550 ;
        RECT 2.065 0.715 2.715 0.905 ;
        RECT 4.035 0.885 4.295 1.775 ;
        RECT 0.975 0.280 1.845 0.560 ;
        RECT 2.025 0.085 2.205 0.545 ;
        RECT 2.460 0.255 2.715 0.715 ;
        RECT 3.520 0.715 4.295 0.885 ;
        RECT 4.515 1.420 4.790 2.135 ;
        RECT 4.960 1.590 5.180 2.465 ;
        RECT 5.430 2.135 6.205 2.465 ;
        RECT 6.445 2.275 6.775 2.635 ;
        RECT 4.515 1.090 4.840 1.420 ;
        RECT 2.940 0.085 3.280 0.555 ;
        RECT 3.520 0.255 3.705 0.715 ;
        RECT 4.515 0.585 4.685 1.090 ;
        RECT 5.010 0.920 5.180 1.590 ;
        RECT 5.605 1.575 5.865 1.955 ;
        RECT 6.035 1.395 6.205 2.135 ;
        RECT 7.100 2.105 7.365 2.450 ;
        RECT 7.655 2.125 8.710 2.635 ;
        RECT 8.880 2.125 9.735 2.460 ;
        RECT 10.045 2.235 10.425 2.635 ;
        RECT 6.425 1.935 7.365 2.105 ;
        RECT 9.565 2.065 9.735 2.125 ;
        RECT 10.645 2.065 10.860 2.450 ;
        RECT 11.135 2.235 11.465 2.635 ;
        RECT 6.425 1.575 6.595 1.935 ;
        RECT 7.190 1.445 7.725 1.765 ;
        RECT 7.910 1.495 8.755 1.955 ;
        RECT 5.485 1.275 6.935 1.395 ;
        RECT 7.950 1.275 8.360 1.325 ;
        RECT 3.930 0.085 4.240 0.545 ;
        RECT 4.460 0.255 4.685 0.585 ;
        RECT 4.855 0.255 5.180 0.920 ;
        RECT 5.400 1.225 8.360 1.275 ;
        RECT 5.400 0.255 5.890 1.225 ;
        RECT 6.060 0.805 6.475 1.015 ;
        RECT 6.750 0.975 8.360 1.225 ;
        RECT 8.535 0.895 8.755 1.495 ;
        RECT 9.115 1.075 9.395 1.905 ;
        RECT 9.565 1.895 11.465 2.065 ;
        RECT 9.685 1.525 11.075 1.725 ;
        RECT 11.245 1.525 11.465 1.895 ;
        RECT 9.685 1.415 9.960 1.525 ;
        RECT 11.685 1.355 11.945 2.465 ;
        RECT 12.170 1.485 12.380 2.635 ;
        RECT 9.610 0.895 9.890 1.245 ;
        RECT 6.060 0.635 7.085 0.805 ;
        RECT 8.535 0.695 9.890 0.895 ;
        RECT 10.140 1.185 11.945 1.355 ;
        RECT 10.140 0.855 10.365 1.185 ;
        RECT 10.605 0.845 11.545 1.015 ;
        RECT 6.060 0.085 6.595 0.465 ;
        RECT 6.775 0.255 7.085 0.635 ;
        RECT 7.540 0.085 8.275 0.690 ;
        RECT 10.605 0.445 10.775 0.845 ;
        RECT 9.160 0.275 10.775 0.445 ;
        RECT 11.220 0.085 11.390 0.545 ;
        RECT 11.765 0.540 11.945 1.185 ;
        RECT 13.160 1.325 13.370 2.465 ;
        RECT 13.725 1.575 13.895 2.635 ;
        RECT 13.160 0.995 14.050 1.325 ;
        RECT 11.560 0.255 11.945 0.540 ;
        RECT 12.170 0.085 12.380 0.885 ;
        RECT 13.160 0.255 13.370 0.995 ;
        RECT 13.690 0.085 13.895 0.825 ;
        RECT 0.000 -0.085 14.720 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 14.405 2.635 14.575 2.805 ;
        RECT 0.630 1.105 0.800 1.275 ;
        RECT 1.675 1.445 1.845 1.615 ;
        RECT 4.125 1.785 4.295 1.955 ;
        RECT 2.645 1.105 2.815 1.275 ;
        RECT 5.010 1.445 5.180 1.615 ;
        RECT 5.605 1.785 5.775 1.955 ;
        RECT 4.585 1.105 4.755 1.275 ;
        RECT 8.205 1.785 8.375 1.955 ;
        RECT 7.445 1.445 7.615 1.615 ;
        RECT 9.735 1.445 9.905 1.615 ;
        RECT 9.225 1.105 9.395 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
        RECT 14.405 -0.085 14.575 0.085 ;
      LAYER met1 ;
        RECT 4.065 1.940 4.405 1.985 ;
        RECT 5.545 1.940 5.885 1.985 ;
        RECT 8.145 1.940 8.435 1.985 ;
        RECT 4.065 1.800 8.435 1.940 ;
        RECT 4.065 1.755 4.405 1.800 ;
        RECT 5.545 1.755 5.885 1.800 ;
        RECT 8.145 1.755 8.435 1.800 ;
        RECT 1.615 1.600 1.955 1.645 ;
        RECT 4.950 1.600 5.240 1.645 ;
        RECT 1.615 1.460 5.240 1.600 ;
        RECT 1.615 1.415 1.955 1.460 ;
        RECT 4.950 1.415 5.240 1.460 ;
        RECT 4.525 1.260 4.815 1.305 ;
        RECT 9.115 1.260 9.455 1.305 ;
        RECT 4.525 1.120 9.455 1.260 ;
        RECT 4.525 1.075 4.815 1.120 ;
        RECT 9.115 1.075 9.455 1.120 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfsbp_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__sdfsbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sdfsbp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.640 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 2.855 1.720 3.335 1.970 ;
        RECT 3.155 1.590 3.335 1.720 ;
        RECT 3.155 1.055 3.815 1.590 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 1.030 0.765 1.425 1.675 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.365 1.675 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.356400 ;
    PORT
      LAYER met1 ;
        RECT 0.570 1.260 0.860 1.305 ;
        RECT 2.585 1.260 2.875 1.305 ;
        RECT 0.570 1.120 2.875 1.260 ;
        RECT 0.570 1.075 0.860 1.120 ;
        RECT 2.585 1.075 2.875 1.120 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277200 ;
    PORT
      LAYER met1 ;
        RECT 7.385 1.600 7.725 1.645 ;
        RECT 9.675 1.600 9.965 1.645 ;
        RECT 7.385 1.460 9.965 1.600 ;
        RECT 7.385 1.415 7.725 1.460 ;
        RECT 9.675 1.415 9.965 1.460 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 15.640 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 7.690 0.785 9.595 1.005 ;
        RECT 12.040 0.785 15.590 1.015 ;
        RECT 0.005 0.105 15.590 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 15.830 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 15.640 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.498000 ;
    PORT
      LAYER li1 ;
        RECT 14.700 1.495 15.080 2.450 ;
        RECT 14.805 0.825 15.080 1.495 ;
        RECT 14.700 0.275 15.080 0.825 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.498000 ;
    PORT
      LAYER li1 ;
        RECT 12.555 0.255 13.000 2.465 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 15.640 2.805 ;
        RECT 0.085 2.025 0.345 2.465 ;
        RECT 0.515 2.195 0.815 2.635 ;
        RECT 1.035 2.255 2.245 2.465 ;
        RECT 1.035 2.025 1.205 2.255 ;
        RECT 2.470 2.085 2.685 2.465 ;
        RECT 2.940 2.140 3.280 2.635 ;
        RECT 0.085 1.845 1.205 2.025 ;
        RECT 1.395 1.870 1.845 2.075 ;
        RECT 0.550 0.765 0.860 1.675 ;
        RECT 0.085 0.085 0.430 0.595 ;
        RECT 1.655 0.560 1.845 1.870 ;
        RECT 2.065 1.770 2.685 2.085 ;
        RECT 3.505 1.955 3.675 2.325 ;
        RECT 3.845 2.275 4.225 2.635 ;
        RECT 4.445 2.135 4.790 2.465 ;
        RECT 3.505 1.775 4.295 1.955 ;
        RECT 2.065 0.905 2.400 1.770 ;
        RECT 2.570 1.075 2.950 1.550 ;
        RECT 2.065 0.715 2.715 0.905 ;
        RECT 4.035 0.885 4.295 1.775 ;
        RECT 0.975 0.280 1.845 0.560 ;
        RECT 2.025 0.085 2.205 0.545 ;
        RECT 2.460 0.255 2.715 0.715 ;
        RECT 3.520 0.715 4.295 0.885 ;
        RECT 4.515 1.420 4.790 2.135 ;
        RECT 4.960 1.590 5.180 2.465 ;
        RECT 5.430 2.135 6.205 2.465 ;
        RECT 6.445 2.275 6.775 2.635 ;
        RECT 4.515 1.090 4.840 1.420 ;
        RECT 2.940 0.085 3.280 0.555 ;
        RECT 3.520 0.255 3.705 0.715 ;
        RECT 4.515 0.585 4.685 1.090 ;
        RECT 5.010 0.920 5.180 1.590 ;
        RECT 5.605 1.575 5.865 1.955 ;
        RECT 6.035 1.395 6.205 2.135 ;
        RECT 7.100 2.105 7.365 2.450 ;
        RECT 7.655 2.125 8.710 2.635 ;
        RECT 8.880 2.125 9.735 2.460 ;
        RECT 10.045 2.235 10.425 2.635 ;
        RECT 6.425 1.935 7.365 2.105 ;
        RECT 9.565 2.065 9.735 2.125 ;
        RECT 10.645 2.065 10.860 2.450 ;
        RECT 11.135 2.235 11.465 2.635 ;
        RECT 6.425 1.575 6.595 1.935 ;
        RECT 7.190 1.445 7.725 1.765 ;
        RECT 7.910 1.495 8.755 1.955 ;
        RECT 5.485 1.275 6.935 1.395 ;
        RECT 7.950 1.275 8.360 1.325 ;
        RECT 3.930 0.085 4.240 0.545 ;
        RECT 4.460 0.255 4.685 0.585 ;
        RECT 4.855 0.255 5.180 0.920 ;
        RECT 5.400 1.225 8.360 1.275 ;
        RECT 5.400 0.255 5.890 1.225 ;
        RECT 6.060 0.805 6.475 1.015 ;
        RECT 6.750 0.975 8.360 1.225 ;
        RECT 8.535 0.895 8.755 1.495 ;
        RECT 9.115 1.075 9.395 1.905 ;
        RECT 9.565 1.895 11.465 2.065 ;
        RECT 9.685 1.525 11.075 1.725 ;
        RECT 11.245 1.525 11.465 1.895 ;
        RECT 9.685 1.415 9.960 1.525 ;
        RECT 11.685 1.355 11.945 2.465 ;
        RECT 12.170 1.485 12.380 2.635 ;
        RECT 13.215 1.485 13.505 2.635 ;
        RECT 9.610 0.895 9.890 1.245 ;
        RECT 6.060 0.635 7.085 0.805 ;
        RECT 8.535 0.695 9.890 0.895 ;
        RECT 10.140 1.185 11.945 1.355 ;
        RECT 10.140 0.855 10.365 1.185 ;
        RECT 10.605 0.845 11.545 1.015 ;
        RECT 6.060 0.085 6.595 0.465 ;
        RECT 6.775 0.255 7.085 0.635 ;
        RECT 7.540 0.085 8.275 0.690 ;
        RECT 10.605 0.445 10.775 0.845 ;
        RECT 9.160 0.275 10.775 0.445 ;
        RECT 11.220 0.085 11.390 0.545 ;
        RECT 11.765 0.540 11.945 1.185 ;
        RECT 13.720 1.325 13.905 2.465 ;
        RECT 14.075 1.635 14.480 2.635 ;
        RECT 15.250 1.485 15.515 2.635 ;
        RECT 13.720 0.995 14.585 1.325 ;
        RECT 11.560 0.255 11.945 0.540 ;
        RECT 12.170 0.085 12.380 0.885 ;
        RECT 13.215 0.085 13.505 0.885 ;
        RECT 13.720 0.255 13.905 0.995 ;
        RECT 14.075 0.085 14.480 0.825 ;
        RECT 15.250 0.085 15.515 0.885 ;
        RECT 0.000 -0.085 15.640 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 14.405 2.635 14.575 2.805 ;
        RECT 14.865 2.635 15.035 2.805 ;
        RECT 15.325 2.635 15.495 2.805 ;
        RECT 0.630 1.105 0.800 1.275 ;
        RECT 1.675 1.445 1.845 1.615 ;
        RECT 4.125 1.785 4.295 1.955 ;
        RECT 2.645 1.105 2.815 1.275 ;
        RECT 5.010 1.445 5.180 1.615 ;
        RECT 5.605 1.785 5.775 1.955 ;
        RECT 4.585 1.105 4.755 1.275 ;
        RECT 8.205 1.785 8.375 1.955 ;
        RECT 7.445 1.445 7.615 1.615 ;
        RECT 9.735 1.445 9.905 1.615 ;
        RECT 9.225 1.105 9.395 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
        RECT 14.405 -0.085 14.575 0.085 ;
        RECT 14.865 -0.085 15.035 0.085 ;
        RECT 15.325 -0.085 15.495 0.085 ;
      LAYER met1 ;
        RECT 4.065 1.940 4.405 1.985 ;
        RECT 5.545 1.940 5.885 1.985 ;
        RECT 8.145 1.940 8.435 1.985 ;
        RECT 4.065 1.800 8.435 1.940 ;
        RECT 4.065 1.755 4.405 1.800 ;
        RECT 5.545 1.755 5.885 1.800 ;
        RECT 8.145 1.755 8.435 1.800 ;
        RECT 1.615 1.600 1.955 1.645 ;
        RECT 4.950 1.600 5.240 1.645 ;
        RECT 1.615 1.460 5.240 1.600 ;
        RECT 1.615 1.415 1.955 1.460 ;
        RECT 4.950 1.415 5.240 1.460 ;
        RECT 4.525 1.260 4.815 1.305 ;
        RECT 9.115 1.260 9.455 1.305 ;
        RECT 4.525 1.120 9.455 1.260 ;
        RECT 4.525 1.075 4.815 1.120 ;
        RECT 9.115 1.075 9.455 1.120 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfsbp_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__sdfstp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sdfstp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.340 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 3.155 1.055 3.815 1.650 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 1.040 0.765 1.485 1.675 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.340 1.675 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.356400 ;
    PORT
      LAYER met1 ;
        RECT 0.580 1.260 0.870 1.305 ;
        RECT 2.585 1.260 2.875 1.305 ;
        RECT 0.580 1.120 2.875 1.260 ;
        RECT 0.580 1.075 0.870 1.120 ;
        RECT 2.585 1.075 2.875 1.120 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277200 ;
    PORT
      LAYER met1 ;
        RECT 7.375 1.600 7.715 1.645 ;
        RECT 9.565 1.600 9.905 1.645 ;
        RECT 7.375 1.460 9.905 1.600 ;
        RECT 7.375 1.415 7.715 1.460 ;
        RECT 9.565 1.415 9.905 1.460 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 13.340 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 7.640 0.785 9.545 1.005 ;
        RECT 12.310 0.785 13.280 1.015 ;
        RECT 0.005 0.105 13.280 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 13.530 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 13.340 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 12.915 0.275 13.240 2.450 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 13.340 2.805 ;
        RECT 0.085 2.025 0.345 2.465 ;
        RECT 0.515 2.195 0.835 2.635 ;
        RECT 1.055 2.255 2.245 2.465 ;
        RECT 1.055 2.025 1.225 2.255 ;
        RECT 2.470 2.085 2.720 2.465 ;
        RECT 2.940 2.140 3.235 2.635 ;
        RECT 0.085 1.845 1.225 2.025 ;
        RECT 1.395 1.845 1.845 2.085 ;
        RECT 0.540 0.765 0.870 1.675 ;
        RECT 1.655 0.595 1.845 1.845 ;
        RECT 2.065 1.770 2.720 2.085 ;
        RECT 3.505 2.000 3.675 2.325 ;
        RECT 3.845 2.275 4.225 2.635 ;
        RECT 4.445 2.135 4.790 2.465 ;
        RECT 3.505 1.830 4.295 2.000 ;
        RECT 2.065 0.905 2.400 1.770 ;
        RECT 2.570 1.075 2.950 1.600 ;
        RECT 2.065 0.715 2.720 0.905 ;
        RECT 4.035 0.885 4.295 1.830 ;
        RECT 0.085 0.085 0.750 0.595 ;
        RECT 0.920 0.255 1.845 0.595 ;
        RECT 2.025 0.085 2.290 0.545 ;
        RECT 2.460 0.255 2.720 0.715 ;
        RECT 3.520 0.715 4.295 0.885 ;
        RECT 4.475 1.420 4.790 2.135 ;
        RECT 4.965 1.590 5.180 2.465 ;
        RECT 5.435 2.135 6.205 2.465 ;
        RECT 6.445 2.275 6.830 2.635 ;
        RECT 4.475 1.085 4.840 1.420 ;
        RECT 2.940 0.085 3.350 0.555 ;
        RECT 3.520 0.255 3.705 0.715 ;
        RECT 3.925 0.085 4.255 0.545 ;
        RECT 4.475 0.255 4.685 1.085 ;
        RECT 5.010 0.780 5.180 1.590 ;
        RECT 5.605 1.575 5.865 1.955 ;
        RECT 6.035 1.395 6.205 2.135 ;
        RECT 7.155 2.105 7.420 2.450 ;
        RECT 7.710 2.125 8.625 2.635 ;
        RECT 8.795 2.125 9.690 2.460 ;
        RECT 9.860 2.235 10.190 2.635 ;
        RECT 6.425 1.935 7.420 2.105 ;
        RECT 9.520 2.065 9.690 2.125 ;
        RECT 10.395 2.065 10.595 2.450 ;
        RECT 10.875 2.235 11.255 2.635 ;
        RECT 6.425 1.575 6.595 1.935 ;
        RECT 7.190 1.445 7.715 1.765 ;
        RECT 7.885 1.670 8.785 1.955 ;
        RECT 4.855 0.255 5.180 0.780 ;
        RECT 5.465 1.275 6.975 1.395 ;
        RECT 7.905 1.275 8.315 1.325 ;
        RECT 5.465 1.225 8.315 1.275 ;
        RECT 5.465 0.255 5.890 1.225 ;
        RECT 6.095 0.805 6.475 1.015 ;
        RECT 6.805 0.975 8.315 1.225 ;
        RECT 8.485 0.905 8.785 1.670 ;
        RECT 8.955 1.075 9.290 1.905 ;
        RECT 9.520 1.895 11.255 2.065 ;
        RECT 9.580 1.545 10.695 1.725 ;
        RECT 10.875 1.605 11.255 1.895 ;
        RECT 9.580 1.425 9.860 1.545 ;
        RECT 11.425 1.365 11.685 2.465 ;
        RECT 9.520 0.905 9.850 1.255 ;
        RECT 6.095 0.635 7.035 0.805 ;
        RECT 6.060 0.085 6.595 0.465 ;
        RECT 6.785 0.255 7.035 0.635 ;
        RECT 7.255 0.085 8.315 0.805 ;
        RECT 8.485 0.720 9.850 0.905 ;
        RECT 10.035 1.195 11.685 1.365 ;
        RECT 10.035 0.855 10.280 1.195 ;
        RECT 10.450 0.785 11.285 1.015 ;
        RECT 10.450 0.545 10.650 0.785 ;
        RECT 11.455 0.585 11.685 1.195 ;
        RECT 9.025 0.275 10.650 0.545 ;
        RECT 10.835 0.085 11.085 0.545 ;
        RECT 11.345 0.255 11.685 0.585 ;
        RECT 11.855 1.325 12.195 2.465 ;
        RECT 12.435 1.845 12.690 2.635 ;
        RECT 11.855 0.995 12.745 1.325 ;
        RECT 11.855 0.255 12.115 0.995 ;
        RECT 12.285 0.085 12.690 0.550 ;
        RECT 0.000 -0.085 13.340 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 0.640 1.105 0.810 1.275 ;
        RECT 1.675 1.445 1.845 1.615 ;
        RECT 4.125 1.785 4.295 1.955 ;
        RECT 2.645 1.105 2.815 1.275 ;
        RECT 5.010 1.445 5.180 1.615 ;
        RECT 5.605 1.785 5.775 1.955 ;
        RECT 4.635 1.100 4.805 1.270 ;
        RECT 8.210 1.785 8.380 1.955 ;
        RECT 7.435 1.445 7.605 1.615 ;
        RECT 9.625 1.445 9.795 1.615 ;
        RECT 9.050 1.105 9.220 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
      LAYER met1 ;
        RECT 4.065 1.940 4.405 1.985 ;
        RECT 5.545 1.940 5.885 1.985 ;
        RECT 8.150 1.940 8.490 1.985 ;
        RECT 4.065 1.800 8.490 1.940 ;
        RECT 4.065 1.755 4.405 1.800 ;
        RECT 5.545 1.755 5.885 1.800 ;
        RECT 8.150 1.755 8.490 1.800 ;
        RECT 1.615 1.600 1.955 1.645 ;
        RECT 4.950 1.600 5.240 1.645 ;
        RECT 1.615 1.460 5.240 1.600 ;
        RECT 1.615 1.415 1.955 1.460 ;
        RECT 4.950 1.415 5.240 1.460 ;
        RECT 4.575 1.260 4.865 1.300 ;
        RECT 8.940 1.260 9.330 1.305 ;
        RECT 4.575 1.120 9.330 1.260 ;
        RECT 4.575 1.070 4.865 1.120 ;
        RECT 8.940 1.075 9.330 1.120 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfstp_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__sdfstp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sdfstp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.260 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 3.155 1.055 3.815 1.650 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 1.040 0.765 1.485 1.675 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.340 1.675 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.356400 ;
    PORT
      LAYER met1 ;
        RECT 0.580 1.260 0.870 1.305 ;
        RECT 2.585 1.260 2.875 1.305 ;
        RECT 0.580 1.120 2.875 1.260 ;
        RECT 0.580 1.075 0.870 1.120 ;
        RECT 2.585 1.075 2.875 1.120 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277200 ;
    PORT
      LAYER met1 ;
        RECT 7.375 1.600 7.715 1.645 ;
        RECT 9.730 1.600 10.070 1.645 ;
        RECT 7.375 1.460 10.070 1.600 ;
        RECT 7.375 1.415 7.715 1.460 ;
        RECT 9.730 1.415 10.070 1.460 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 14.260 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 7.690 0.785 9.695 1.005 ;
        RECT 12.640 0.785 14.175 1.015 ;
        RECT 0.005 0.105 14.175 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 14.450 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 14.260 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.498000 ;
    PORT
      LAYER li1 ;
        RECT 13.245 1.495 13.655 2.450 ;
        RECT 13.350 0.825 13.655 1.495 ;
        RECT 13.245 0.275 13.655 0.825 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 14.260 2.805 ;
        RECT 0.085 2.025 0.345 2.465 ;
        RECT 0.515 2.195 0.835 2.635 ;
        RECT 1.055 2.255 2.245 2.465 ;
        RECT 1.055 2.025 1.225 2.255 ;
        RECT 2.470 2.085 2.720 2.465 ;
        RECT 2.940 2.140 3.235 2.635 ;
        RECT 0.085 1.845 1.225 2.025 ;
        RECT 1.395 1.845 1.845 2.085 ;
        RECT 0.540 0.765 0.870 1.675 ;
        RECT 1.655 0.595 1.845 1.845 ;
        RECT 2.065 1.770 2.720 2.085 ;
        RECT 3.505 2.000 3.675 2.325 ;
        RECT 3.845 2.275 4.225 2.635 ;
        RECT 4.445 2.135 4.790 2.465 ;
        RECT 3.505 1.830 4.295 2.000 ;
        RECT 2.065 0.905 2.400 1.770 ;
        RECT 2.570 1.075 2.950 1.600 ;
        RECT 2.065 0.715 2.720 0.905 ;
        RECT 4.035 0.885 4.295 1.830 ;
        RECT 0.085 0.085 0.750 0.595 ;
        RECT 0.920 0.255 1.845 0.595 ;
        RECT 2.025 0.085 2.290 0.545 ;
        RECT 2.460 0.255 2.720 0.715 ;
        RECT 3.520 0.715 4.295 0.885 ;
        RECT 4.475 1.420 4.790 2.135 ;
        RECT 4.965 1.590 5.180 2.465 ;
        RECT 5.435 2.135 6.205 2.465 ;
        RECT 6.445 2.275 6.830 2.635 ;
        RECT 4.475 1.085 4.840 1.420 ;
        RECT 2.940 0.085 3.350 0.555 ;
        RECT 3.520 0.255 3.705 0.715 ;
        RECT 3.925 0.085 4.255 0.545 ;
        RECT 4.475 0.255 4.685 1.085 ;
        RECT 5.010 0.780 5.180 1.590 ;
        RECT 5.605 1.575 5.865 1.955 ;
        RECT 6.035 1.395 6.205 2.135 ;
        RECT 7.155 2.105 7.420 2.450 ;
        RECT 7.710 2.125 8.765 2.635 ;
        RECT 8.935 2.125 9.840 2.460 ;
        RECT 10.060 2.235 10.440 2.635 ;
        RECT 6.425 1.935 7.420 2.105 ;
        RECT 9.670 2.065 9.840 2.125 ;
        RECT 10.610 2.065 11.015 2.450 ;
        RECT 11.205 2.235 11.585 2.635 ;
        RECT 6.425 1.575 6.595 1.935 ;
        RECT 7.190 1.445 7.715 1.765 ;
        RECT 7.885 1.670 8.885 1.955 ;
        RECT 4.855 0.255 5.180 0.780 ;
        RECT 5.465 1.275 6.975 1.395 ;
        RECT 8.005 1.275 8.415 1.325 ;
        RECT 5.465 1.225 8.415 1.275 ;
        RECT 5.465 0.255 5.890 1.225 ;
        RECT 6.095 0.805 6.475 1.015 ;
        RECT 6.805 0.975 8.415 1.225 ;
        RECT 8.585 0.905 8.885 1.670 ;
        RECT 9.175 1.075 9.500 1.905 ;
        RECT 9.670 1.895 11.585 2.065 ;
        RECT 9.730 1.545 10.995 1.725 ;
        RECT 11.205 1.605 11.585 1.895 ;
        RECT 9.730 1.425 10.035 1.545 ;
        RECT 11.755 1.365 12.015 2.465 ;
        RECT 9.670 0.905 10.005 1.255 ;
        RECT 6.095 0.635 7.035 0.805 ;
        RECT 6.060 0.085 6.595 0.465 ;
        RECT 6.785 0.255 7.035 0.635 ;
        RECT 7.255 0.085 8.415 0.805 ;
        RECT 8.585 0.720 10.005 0.905 ;
        RECT 10.220 1.195 12.015 1.365 ;
        RECT 10.220 0.855 10.480 1.195 ;
        RECT 10.710 0.785 11.615 1.015 ;
        RECT 10.710 0.545 10.910 0.785 ;
        RECT 11.785 0.585 12.015 1.195 ;
        RECT 9.265 0.275 10.910 0.545 ;
        RECT 11.165 0.085 11.415 0.545 ;
        RECT 11.675 0.255 12.015 0.585 ;
        RECT 12.185 1.325 12.525 2.465 ;
        RECT 12.765 1.845 13.020 2.635 ;
        RECT 13.825 1.495 13.995 2.635 ;
        RECT 12.185 0.995 13.125 1.325 ;
        RECT 12.185 0.255 12.445 0.995 ;
        RECT 12.615 0.085 13.020 0.550 ;
        RECT 13.825 0.085 13.995 0.885 ;
        RECT 0.000 -0.085 14.260 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 0.640 1.105 0.810 1.275 ;
        RECT 1.675 1.445 1.845 1.615 ;
        RECT 4.125 1.785 4.295 1.955 ;
        RECT 2.645 1.105 2.815 1.275 ;
        RECT 5.010 1.445 5.180 1.615 ;
        RECT 5.605 1.785 5.775 1.955 ;
        RECT 4.635 1.100 4.805 1.270 ;
        RECT 8.210 1.785 8.380 1.955 ;
        RECT 7.435 1.445 7.605 1.615 ;
        RECT 9.790 1.445 9.960 1.615 ;
        RECT 9.280 1.105 9.450 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
      LAYER met1 ;
        RECT 4.065 1.940 4.405 1.985 ;
        RECT 5.545 1.940 5.885 1.985 ;
        RECT 8.150 1.940 8.490 1.985 ;
        RECT 4.065 1.800 8.490 1.940 ;
        RECT 4.065 1.755 4.405 1.800 ;
        RECT 5.545 1.755 5.885 1.800 ;
        RECT 8.150 1.755 8.490 1.800 ;
        RECT 1.615 1.600 1.955 1.645 ;
        RECT 4.950 1.600 5.240 1.645 ;
        RECT 1.615 1.460 5.240 1.600 ;
        RECT 1.615 1.415 1.955 1.460 ;
        RECT 4.950 1.415 5.240 1.460 ;
        RECT 4.575 1.260 4.865 1.300 ;
        RECT 9.170 1.260 9.560 1.305 ;
        RECT 4.575 1.120 9.560 1.260 ;
        RECT 4.575 1.070 4.865 1.120 ;
        RECT 9.170 1.075 9.560 1.120 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfstp_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__sdfstp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sdfstp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.180 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 3.155 1.055 3.815 1.650 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 1.040 0.765 1.485 1.675 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.340 1.675 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.356400 ;
    PORT
      LAYER met1 ;
        RECT 0.580 1.260 0.870 1.305 ;
        RECT 2.585 1.260 2.875 1.305 ;
        RECT 0.580 1.120 2.875 1.260 ;
        RECT 0.580 1.075 0.870 1.120 ;
        RECT 2.585 1.075 2.875 1.120 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277200 ;
    PORT
      LAYER met1 ;
        RECT 7.375 1.600 7.715 1.645 ;
        RECT 9.730 1.600 10.070 1.645 ;
        RECT 7.375 1.460 10.070 1.600 ;
        RECT 7.375 1.415 7.715 1.460 ;
        RECT 9.730 1.415 10.070 1.460 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 15.180 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 7.690 0.785 9.695 1.005 ;
        RECT 12.105 0.785 15.120 1.015 ;
        RECT 0.005 0.105 15.120 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 15.370 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 15.180 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.996000 ;
    PORT
      LAYER li1 ;
        RECT 13.240 1.495 13.570 2.450 ;
        RECT 13.345 1.325 13.570 1.495 ;
        RECT 14.130 1.325 14.610 2.465 ;
        RECT 13.345 1.055 14.610 1.325 ;
        RECT 13.345 0.825 13.570 1.055 ;
        RECT 13.240 0.275 13.570 0.825 ;
        RECT 14.130 0.255 14.610 1.055 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 15.180 2.805 ;
        RECT 0.085 2.025 0.345 2.465 ;
        RECT 0.515 2.195 0.835 2.635 ;
        RECT 1.055 2.255 2.245 2.465 ;
        RECT 1.055 2.025 1.225 2.255 ;
        RECT 2.470 2.085 2.720 2.465 ;
        RECT 2.940 2.140 3.235 2.635 ;
        RECT 0.085 1.845 1.225 2.025 ;
        RECT 1.395 1.845 1.845 2.085 ;
        RECT 0.540 0.765 0.870 1.675 ;
        RECT 1.655 0.595 1.845 1.845 ;
        RECT 2.065 1.770 2.720 2.085 ;
        RECT 3.505 2.000 3.675 2.325 ;
        RECT 3.845 2.275 4.225 2.635 ;
        RECT 4.445 2.135 4.790 2.465 ;
        RECT 3.505 1.830 4.295 2.000 ;
        RECT 2.065 0.905 2.400 1.770 ;
        RECT 2.570 1.075 2.950 1.600 ;
        RECT 2.065 0.715 2.720 0.905 ;
        RECT 4.035 0.885 4.295 1.830 ;
        RECT 0.085 0.085 0.750 0.595 ;
        RECT 0.920 0.255 1.845 0.595 ;
        RECT 2.025 0.085 2.290 0.545 ;
        RECT 2.460 0.255 2.720 0.715 ;
        RECT 3.520 0.715 4.295 0.885 ;
        RECT 4.475 1.420 4.790 2.135 ;
        RECT 4.965 1.590 5.180 2.465 ;
        RECT 5.435 2.135 6.205 2.465 ;
        RECT 6.445 2.275 6.830 2.635 ;
        RECT 4.475 1.085 4.840 1.420 ;
        RECT 2.940 0.085 3.350 0.555 ;
        RECT 3.520 0.255 3.705 0.715 ;
        RECT 3.925 0.085 4.255 0.545 ;
        RECT 4.475 0.255 4.685 1.085 ;
        RECT 5.010 0.780 5.180 1.590 ;
        RECT 5.605 1.575 5.865 1.955 ;
        RECT 6.035 1.395 6.205 2.135 ;
        RECT 7.155 2.105 7.420 2.450 ;
        RECT 7.710 2.125 8.765 2.635 ;
        RECT 8.935 2.125 9.840 2.460 ;
        RECT 10.060 2.235 10.440 2.635 ;
        RECT 6.425 1.935 7.420 2.105 ;
        RECT 9.670 2.065 9.840 2.125 ;
        RECT 10.610 2.065 11.015 2.450 ;
        RECT 11.205 2.235 11.585 2.635 ;
        RECT 6.425 1.575 6.595 1.935 ;
        RECT 7.190 1.445 7.715 1.765 ;
        RECT 7.885 1.670 8.885 1.955 ;
        RECT 4.855 0.255 5.180 0.780 ;
        RECT 5.465 1.275 6.975 1.395 ;
        RECT 8.005 1.275 8.415 1.325 ;
        RECT 5.465 1.225 8.415 1.275 ;
        RECT 5.465 0.255 5.890 1.225 ;
        RECT 6.095 0.805 6.475 1.015 ;
        RECT 6.805 0.975 8.415 1.225 ;
        RECT 8.585 0.905 8.885 1.670 ;
        RECT 9.175 1.075 9.500 1.905 ;
        RECT 9.670 1.895 11.585 2.065 ;
        RECT 9.730 1.545 10.995 1.725 ;
        RECT 11.205 1.605 11.585 1.895 ;
        RECT 9.730 1.425 10.035 1.545 ;
        RECT 11.755 1.365 12.015 2.465 ;
        RECT 9.670 0.905 10.005 1.255 ;
        RECT 6.095 0.635 7.035 0.805 ;
        RECT 6.060 0.085 6.595 0.465 ;
        RECT 6.785 0.255 7.035 0.635 ;
        RECT 7.255 0.085 8.415 0.805 ;
        RECT 8.585 0.720 10.005 0.905 ;
        RECT 10.220 1.195 12.015 1.365 ;
        RECT 10.220 0.855 10.480 1.195 ;
        RECT 10.710 0.785 11.615 1.015 ;
        RECT 10.710 0.545 10.910 0.785 ;
        RECT 11.785 0.585 12.015 1.195 ;
        RECT 9.265 0.275 10.910 0.545 ;
        RECT 11.165 0.085 11.415 0.545 ;
        RECT 11.675 0.255 12.015 0.585 ;
        RECT 12.185 1.325 12.445 2.465 ;
        RECT 12.615 1.495 13.020 2.635 ;
        RECT 13.790 1.495 13.960 2.635 ;
        RECT 14.780 1.495 15.065 2.635 ;
        RECT 12.185 0.995 13.125 1.325 ;
        RECT 12.185 0.255 12.445 0.995 ;
        RECT 12.615 0.085 13.020 0.825 ;
        RECT 13.790 0.085 13.960 0.885 ;
        RECT 14.780 0.085 15.065 0.885 ;
        RECT 0.000 -0.085 15.180 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 14.405 2.635 14.575 2.805 ;
        RECT 14.865 2.635 15.035 2.805 ;
        RECT 0.640 1.105 0.810 1.275 ;
        RECT 1.675 1.445 1.845 1.615 ;
        RECT 4.125 1.785 4.295 1.955 ;
        RECT 2.645 1.105 2.815 1.275 ;
        RECT 5.010 1.445 5.180 1.615 ;
        RECT 5.605 1.785 5.775 1.955 ;
        RECT 4.635 1.100 4.805 1.270 ;
        RECT 8.210 1.785 8.380 1.955 ;
        RECT 7.435 1.445 7.605 1.615 ;
        RECT 9.790 1.445 9.960 1.615 ;
        RECT 9.280 1.105 9.450 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
        RECT 14.405 -0.085 14.575 0.085 ;
        RECT 14.865 -0.085 15.035 0.085 ;
      LAYER met1 ;
        RECT 4.065 1.940 4.405 1.985 ;
        RECT 5.545 1.940 5.885 1.985 ;
        RECT 8.150 1.940 8.490 1.985 ;
        RECT 4.065 1.800 8.490 1.940 ;
        RECT 4.065 1.755 4.405 1.800 ;
        RECT 5.545 1.755 5.885 1.800 ;
        RECT 8.150 1.755 8.490 1.800 ;
        RECT 1.615 1.600 1.955 1.645 ;
        RECT 4.950 1.600 5.240 1.645 ;
        RECT 1.615 1.460 5.240 1.600 ;
        RECT 1.615 1.415 1.955 1.460 ;
        RECT 4.950 1.415 5.240 1.460 ;
        RECT 4.575 1.260 4.865 1.300 ;
        RECT 9.170 1.260 9.560 1.305 ;
        RECT 4.575 1.120 9.560 1.260 ;
        RECT 4.575 1.070 4.865 1.120 ;
        RECT 9.170 1.075 9.560 1.120 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfstp_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__sdfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sdfxbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.960 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 2.755 1.355 3.125 1.685 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 3.815 1.055 4.345 1.655 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.356400 ;
    PORT
      LAYER li1 ;
        RECT 1.860 0.785 2.030 1.685 ;
        RECT 3.315 0.785 3.535 1.115 ;
        RECT 1.860 0.615 3.535 0.785 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.960 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 6.325 0.785 7.285 1.005 ;
        RECT 8.980 0.785 11.955 1.015 ;
        RECT 0.005 0.725 4.435 0.785 ;
        RECT 5.545 0.725 11.955 0.785 ;
        RECT 0.005 0.105 11.955 0.725 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 12.150 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.960 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 9.980 1.505 10.440 2.465 ;
        RECT 10.220 0.825 10.440 1.505 ;
        RECT 9.960 0.305 10.440 0.825 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 11.615 0.265 11.870 2.325 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 11.960 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.895 2.635 ;
        RECT 0.175 1.795 0.895 1.965 ;
        RECT 0.665 0.970 0.895 1.795 ;
        RECT 0.665 0.805 0.860 0.970 ;
        RECT 0.175 0.635 0.860 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.115 0.345 1.285 2.465 ;
        RECT 1.520 2.075 1.805 2.445 ;
        RECT 1.975 2.245 2.355 2.635 ;
        RECT 2.875 2.245 3.870 2.415 ;
        RECT 1.520 1.860 3.530 2.075 ;
        RECT 1.520 0.445 1.690 1.860 ;
        RECT 2.250 1.125 2.420 1.860 ;
        RECT 3.335 1.685 3.530 1.860 ;
        RECT 3.700 1.995 3.870 2.245 ;
        RECT 4.090 2.165 4.260 2.635 ;
        RECT 4.515 2.070 4.800 2.440 ;
        RECT 4.995 2.190 6.215 2.360 ;
        RECT 4.515 1.995 4.685 2.070 ;
        RECT 3.700 1.825 4.685 1.995 ;
        RECT 3.335 1.355 3.555 1.685 ;
        RECT 2.250 0.955 2.695 1.125 ;
        RECT 4.515 0.885 4.685 1.825 ;
        RECT 3.705 0.715 4.685 0.885 ;
        RECT 3.705 0.445 3.875 0.715 ;
        RECT 1.520 0.255 1.905 0.445 ;
        RECT 2.145 0.085 2.475 0.445 ;
        RECT 3.050 0.275 3.875 0.445 ;
        RECT 4.095 0.085 4.295 0.545 ;
        RECT 4.515 0.535 4.685 0.715 ;
        RECT 4.855 1.035 5.145 1.905 ;
        RECT 5.335 1.655 5.825 2.010 ;
        RECT 5.995 1.575 6.215 2.190 ;
        RECT 6.385 1.835 6.555 2.635 ;
        RECT 6.725 2.135 7.025 2.465 ;
        RECT 7.250 2.165 8.285 2.335 ;
        RECT 5.995 1.485 6.555 1.575 ;
        RECT 5.705 1.315 6.555 1.485 ;
        RECT 4.855 0.705 5.485 1.035 ;
        RECT 5.705 0.535 5.875 1.315 ;
        RECT 6.385 1.245 6.555 1.315 ;
        RECT 6.095 1.065 6.265 1.095 ;
        RECT 6.725 1.065 6.945 2.135 ;
        RECT 7.115 1.245 7.355 1.965 ;
        RECT 7.525 1.575 7.895 1.905 ;
        RECT 6.095 0.765 6.945 1.065 ;
        RECT 7.525 1.035 7.715 1.575 ;
        RECT 8.115 1.405 8.285 2.165 ;
        RECT 8.515 2.135 8.820 2.635 ;
        RECT 9.110 1.905 9.400 2.455 ;
        RECT 8.485 1.575 9.400 1.905 ;
        RECT 9.620 1.625 9.790 2.635 ;
        RECT 4.515 0.365 4.865 0.535 ;
        RECT 5.085 0.365 5.875 0.535 ;
        RECT 6.175 0.085 6.545 0.585 ;
        RECT 6.725 0.535 6.945 0.765 ;
        RECT 7.115 0.705 7.715 1.035 ;
        RECT 7.935 1.325 8.285 1.405 ;
        RECT 9.215 1.325 9.400 1.575 ;
        RECT 10.610 1.325 10.860 2.425 ;
        RECT 11.090 1.495 11.395 2.635 ;
        RECT 7.935 0.995 9.045 1.325 ;
        RECT 9.215 0.995 10.050 1.325 ;
        RECT 10.610 0.995 11.440 1.325 ;
        RECT 7.935 0.535 8.155 0.995 ;
        RECT 9.215 0.825 9.400 0.995 ;
        RECT 6.725 0.365 7.235 0.535 ;
        RECT 7.515 0.365 8.155 0.535 ;
        RECT 8.380 0.085 8.800 0.615 ;
        RECT 9.070 0.300 9.400 0.825 ;
        RECT 9.620 0.085 9.790 0.695 ;
        RECT 10.610 0.345 10.860 0.995 ;
        RECT 11.065 0.085 11.395 0.805 ;
        RECT 0.000 -0.085 11.960 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 0.695 1.785 0.865 1.955 ;
        RECT 1.115 0.425 1.285 0.595 ;
        RECT 5.615 1.785 5.785 1.955 ;
        RECT 5.205 0.765 5.375 0.935 ;
        RECT 7.175 1.785 7.345 1.955 ;
        RECT 7.185 0.765 7.355 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
      LAYER met1 ;
        RECT 0.635 1.940 0.925 1.985 ;
        RECT 5.555 1.940 5.845 1.985 ;
        RECT 7.115 1.940 7.405 1.985 ;
        RECT 0.635 1.800 7.405 1.940 ;
        RECT 0.635 1.755 0.925 1.800 ;
        RECT 5.555 1.755 5.845 1.800 ;
        RECT 7.115 1.755 7.405 1.800 ;
        RECT 5.145 0.920 5.435 0.965 ;
        RECT 7.125 0.920 7.415 0.965 ;
        RECT 5.145 0.780 7.415 0.920 ;
        RECT 5.145 0.735 5.435 0.780 ;
        RECT 7.125 0.735 7.415 0.780 ;
        RECT 1.005 0.580 1.345 0.625 ;
        RECT 5.145 0.580 5.285 0.735 ;
        RECT 1.005 0.440 5.285 0.580 ;
        RECT 1.005 0.395 1.345 0.440 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfxbp_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__sdfxbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sdfxbp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.340 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 2.755 1.355 3.125 1.685 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 3.815 1.055 4.345 1.655 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.356400 ;
    PORT
      LAYER li1 ;
        RECT 1.860 0.785 2.030 1.685 ;
        RECT 3.315 0.785 3.535 1.115 ;
        RECT 1.860 0.615 3.535 0.785 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 13.340 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 6.325 0.785 7.285 1.005 ;
        RECT 8.980 0.785 13.325 1.015 ;
        RECT 0.005 0.725 4.435 0.785 ;
        RECT 5.545 0.725 13.325 0.785 ;
        RECT 0.005 0.105 13.325 0.725 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 13.530 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 13.340 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.498000 ;
    PORT
      LAYER li1 ;
        RECT 10.210 0.255 10.490 2.455 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.498000 ;
    PORT
      LAYER li1 ;
        RECT 12.515 0.265 12.785 2.325 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 13.340 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.895 2.635 ;
        RECT 0.175 1.795 0.895 1.965 ;
        RECT 0.665 0.970 0.895 1.795 ;
        RECT 0.665 0.805 0.860 0.970 ;
        RECT 0.175 0.635 0.860 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.115 0.345 1.285 2.465 ;
        RECT 1.520 2.075 1.805 2.445 ;
        RECT 1.975 2.245 2.355 2.635 ;
        RECT 2.875 2.245 3.870 2.415 ;
        RECT 1.520 1.860 3.530 2.075 ;
        RECT 1.520 0.445 1.690 1.860 ;
        RECT 2.250 1.125 2.420 1.860 ;
        RECT 3.335 1.685 3.530 1.860 ;
        RECT 3.700 1.995 3.870 2.245 ;
        RECT 4.090 2.165 4.260 2.635 ;
        RECT 4.515 2.070 4.800 2.440 ;
        RECT 4.995 2.190 6.215 2.360 ;
        RECT 4.515 1.995 4.685 2.070 ;
        RECT 3.700 1.825 4.685 1.995 ;
        RECT 3.335 1.355 3.555 1.685 ;
        RECT 2.250 0.955 2.695 1.125 ;
        RECT 4.515 0.885 4.685 1.825 ;
        RECT 3.705 0.715 4.685 0.885 ;
        RECT 3.705 0.445 3.875 0.715 ;
        RECT 1.520 0.255 1.905 0.445 ;
        RECT 2.145 0.085 2.475 0.445 ;
        RECT 3.050 0.275 3.875 0.445 ;
        RECT 4.095 0.085 4.295 0.545 ;
        RECT 4.515 0.535 4.685 0.715 ;
        RECT 4.855 1.035 5.145 1.905 ;
        RECT 5.335 1.655 5.825 2.010 ;
        RECT 5.995 1.575 6.215 2.190 ;
        RECT 6.385 1.835 6.555 2.635 ;
        RECT 6.725 2.135 7.025 2.465 ;
        RECT 7.250 2.165 8.285 2.335 ;
        RECT 5.995 1.485 6.555 1.575 ;
        RECT 5.705 1.315 6.555 1.485 ;
        RECT 4.855 0.705 5.485 1.035 ;
        RECT 5.705 0.535 5.875 1.315 ;
        RECT 6.385 1.245 6.555 1.315 ;
        RECT 6.095 1.065 6.265 1.095 ;
        RECT 6.725 1.065 6.945 2.135 ;
        RECT 7.115 1.245 7.355 1.965 ;
        RECT 7.525 1.575 7.895 1.905 ;
        RECT 6.095 0.765 6.945 1.065 ;
        RECT 7.525 1.035 7.715 1.575 ;
        RECT 8.115 1.405 8.285 2.165 ;
        RECT 8.515 2.135 8.820 2.635 ;
        RECT 9.070 1.905 9.400 2.455 ;
        RECT 8.485 1.575 9.400 1.905 ;
        RECT 9.570 1.625 9.990 2.635 ;
        RECT 10.690 1.615 10.860 2.635 ;
        RECT 4.515 0.365 4.865 0.535 ;
        RECT 5.085 0.365 5.875 0.535 ;
        RECT 6.175 0.085 6.545 0.585 ;
        RECT 6.725 0.535 6.945 0.765 ;
        RECT 7.115 0.705 7.715 1.035 ;
        RECT 7.935 1.325 8.285 1.405 ;
        RECT 9.215 1.325 9.400 1.575 ;
        RECT 11.130 1.325 11.460 2.425 ;
        RECT 11.690 1.495 12.295 2.635 ;
        RECT 12.985 1.395 13.155 2.635 ;
        RECT 7.935 0.995 9.045 1.325 ;
        RECT 9.215 0.995 10.000 1.325 ;
        RECT 11.130 0.995 12.340 1.325 ;
        RECT 7.935 0.535 8.155 0.995 ;
        RECT 9.215 0.825 9.400 0.995 ;
        RECT 6.725 0.365 7.235 0.535 ;
        RECT 7.515 0.365 8.155 0.535 ;
        RECT 8.380 0.085 8.800 0.615 ;
        RECT 9.035 0.300 9.400 0.825 ;
        RECT 9.570 0.085 9.990 0.695 ;
        RECT 10.680 0.085 10.910 0.690 ;
        RECT 11.130 0.345 11.380 0.995 ;
        RECT 11.665 0.085 12.295 0.805 ;
        RECT 12.985 0.085 13.155 0.955 ;
        RECT 0.000 -0.085 13.340 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 0.695 1.785 0.865 1.955 ;
        RECT 1.115 0.425 1.285 0.595 ;
        RECT 5.615 1.785 5.785 1.955 ;
        RECT 5.145 0.765 5.315 0.935 ;
        RECT 7.175 1.785 7.345 1.955 ;
        RECT 7.185 0.765 7.355 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
      LAYER met1 ;
        RECT 0.635 1.940 0.925 1.985 ;
        RECT 5.555 1.940 5.845 1.985 ;
        RECT 7.115 1.940 7.405 1.985 ;
        RECT 0.635 1.800 7.405 1.940 ;
        RECT 0.635 1.755 0.925 1.800 ;
        RECT 5.555 1.755 5.845 1.800 ;
        RECT 7.115 1.755 7.405 1.800 ;
        RECT 5.085 0.920 5.375 0.965 ;
        RECT 7.125 0.920 7.415 0.965 ;
        RECT 5.085 0.780 7.415 0.920 ;
        RECT 5.085 0.735 5.375 0.780 ;
        RECT 7.125 0.735 7.415 0.780 ;
        RECT 1.005 0.580 1.345 0.625 ;
        RECT 5.085 0.580 5.225 0.735 ;
        RECT 1.005 0.440 5.225 0.580 ;
        RECT 1.005 0.395 1.345 0.440 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfxbp_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__sdfxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sdfxtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.580 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 2.745 1.355 3.150 1.685 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 3.725 1.035 4.095 1.655 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.356400 ;
    PORT
      LAYER li1 ;
        RECT 1.880 0.785 2.215 1.685 ;
        RECT 3.335 0.785 3.505 1.115 ;
        RECT 1.880 0.615 3.505 0.785 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.580 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 6.275 0.785 7.220 1.005 ;
        RECT 8.950 0.785 10.400 1.015 ;
        RECT 0.005 0.725 4.475 0.785 ;
        RECT 5.565 0.725 10.400 0.785 ;
        RECT 0.005 0.105 10.400 0.725 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.770 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.580 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.471500 ;
    PORT
      LAYER li1 ;
        RECT 9.930 1.545 10.470 2.395 ;
        RECT 10.230 0.820 10.470 1.545 ;
        RECT 9.930 0.305 10.470 0.820 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.580 2.805 ;
        RECT 0.180 1.965 0.350 2.465 ;
        RECT 0.520 2.135 0.900 2.635 ;
        RECT 0.180 1.795 0.895 1.965 ;
        RECT 0.665 0.805 0.895 1.795 ;
        RECT 0.175 0.635 0.895 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.115 0.345 1.345 2.465 ;
        RECT 1.535 2.075 1.810 2.445 ;
        RECT 1.980 2.245 2.360 2.635 ;
        RECT 2.895 2.245 3.890 2.415 ;
        RECT 1.535 1.860 3.540 2.075 ;
        RECT 1.535 0.445 1.705 1.860 ;
        RECT 2.385 1.125 2.555 1.860 ;
        RECT 3.330 1.355 3.540 1.860 ;
        RECT 3.720 1.995 3.890 2.245 ;
        RECT 4.110 2.165 4.280 2.635 ;
        RECT 4.565 2.065 4.800 2.440 ;
        RECT 5.045 2.190 6.230 2.360 ;
        RECT 4.565 1.995 4.735 2.065 ;
        RECT 3.720 1.825 4.735 1.995 ;
        RECT 2.385 0.955 2.715 1.125 ;
        RECT 4.565 0.865 4.735 1.825 ;
        RECT 3.725 0.695 4.735 0.865 ;
        RECT 4.905 1.035 5.195 1.905 ;
        RECT 5.385 1.655 5.875 2.010 ;
        RECT 6.045 1.575 6.230 2.190 ;
        RECT 6.400 1.835 6.570 2.635 ;
        RECT 6.045 1.485 6.685 1.575 ;
        RECT 5.705 1.315 6.685 1.485 ;
        RECT 4.905 0.705 5.535 1.035 ;
        RECT 3.725 0.445 3.895 0.695 ;
        RECT 4.565 0.535 4.735 0.695 ;
        RECT 5.705 0.535 5.875 1.315 ;
        RECT 6.855 1.095 7.060 2.465 ;
        RECT 7.250 2.165 8.285 2.335 ;
        RECT 7.230 1.245 7.470 1.965 ;
        RECT 6.045 0.765 7.060 1.095 ;
        RECT 7.735 1.035 7.945 1.905 ;
        RECT 1.535 0.275 1.905 0.445 ;
        RECT 2.075 0.085 2.405 0.445 ;
        RECT 3.070 0.275 3.895 0.445 ;
        RECT 4.115 0.085 4.315 0.525 ;
        RECT 4.565 0.365 4.915 0.535 ;
        RECT 5.135 0.365 5.875 0.535 ;
        RECT 6.225 0.085 6.595 0.585 ;
        RECT 6.775 0.535 7.060 0.765 ;
        RECT 7.250 0.705 7.945 1.035 ;
        RECT 8.115 1.325 8.285 2.165 ;
        RECT 8.465 2.135 8.770 2.635 ;
        RECT 9.120 1.905 9.405 2.455 ;
        RECT 8.455 1.575 9.405 1.905 ;
        RECT 9.590 1.625 9.760 2.635 ;
        RECT 9.220 1.325 9.405 1.575 ;
        RECT 8.115 0.995 9.050 1.325 ;
        RECT 9.220 0.995 10.030 1.325 ;
        RECT 8.115 0.535 8.285 0.995 ;
        RECT 9.220 0.825 9.400 0.995 ;
        RECT 6.775 0.365 7.260 0.535 ;
        RECT 7.455 0.365 8.285 0.535 ;
        RECT 8.455 0.085 8.770 0.615 ;
        RECT 9.040 0.300 9.400 0.825 ;
        RECT 9.590 0.085 9.760 0.695 ;
        RECT 0.000 -0.085 10.580 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 0.665 1.740 0.835 1.910 ;
        RECT 1.155 0.720 1.325 0.890 ;
        RECT 5.665 1.740 5.835 1.910 ;
        RECT 5.155 0.720 5.325 0.890 ;
        RECT 7.240 1.740 7.410 1.910 ;
        RECT 7.310 0.720 7.480 0.890 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
      LAYER met1 ;
        RECT 0.605 1.800 7.470 1.940 ;
        RECT 0.605 1.710 0.895 1.800 ;
        RECT 5.555 1.710 5.895 1.800 ;
        RECT 7.130 1.710 7.470 1.800 ;
        RECT 1.095 0.780 7.540 0.920 ;
        RECT 1.095 0.690 1.385 0.780 ;
        RECT 5.045 0.690 5.385 0.780 ;
        RECT 7.230 0.690 7.540 0.780 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfxtp_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__sdfxtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sdfxtp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.040 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 2.745 1.355 3.150 1.685 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 3.725 1.035 4.095 1.655 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.356400 ;
    PORT
      LAYER li1 ;
        RECT 1.880 0.785 2.215 1.685 ;
        RECT 3.335 0.785 3.505 1.115 ;
        RECT 1.880 0.615 3.505 0.785 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.040 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 6.375 0.785 7.335 1.005 ;
        RECT 9.050 0.785 11.035 1.015 ;
        RECT 0.005 0.725 4.475 0.785 ;
        RECT 5.595 0.725 11.035 0.785 ;
        RECT 0.005 0.105 11.035 0.725 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 11.230 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.040 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.530500 ;
    PORT
      LAYER li1 ;
        RECT 10.030 1.545 10.500 2.395 ;
        RECT 10.330 0.820 10.500 1.545 ;
        RECT 10.030 0.305 10.500 0.820 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 11.040 2.805 ;
        RECT 0.180 1.965 0.350 2.465 ;
        RECT 0.520 2.135 0.900 2.635 ;
        RECT 0.180 1.795 0.895 1.965 ;
        RECT 0.665 0.805 0.895 1.795 ;
        RECT 0.175 0.635 0.895 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.115 0.345 1.345 2.465 ;
        RECT 1.535 2.075 1.810 2.445 ;
        RECT 1.980 2.245 2.360 2.635 ;
        RECT 2.895 2.245 3.890 2.415 ;
        RECT 1.535 1.860 3.525 2.075 ;
        RECT 1.535 0.445 1.705 1.860 ;
        RECT 2.385 1.125 2.555 1.860 ;
        RECT 3.330 1.355 3.525 1.860 ;
        RECT 3.720 1.995 3.890 2.245 ;
        RECT 4.110 2.165 4.280 2.635 ;
        RECT 4.565 2.065 4.800 2.440 ;
        RECT 5.045 2.190 6.265 2.360 ;
        RECT 4.565 1.995 4.735 2.065 ;
        RECT 3.720 1.825 4.735 1.995 ;
        RECT 2.385 0.955 2.715 1.125 ;
        RECT 4.565 0.865 4.735 1.825 ;
        RECT 3.725 0.695 4.735 0.865 ;
        RECT 4.905 1.035 5.195 1.905 ;
        RECT 5.385 1.655 5.875 2.010 ;
        RECT 6.045 1.575 6.265 2.190 ;
        RECT 6.435 1.835 6.605 2.635 ;
        RECT 6.775 2.135 7.075 2.465 ;
        RECT 7.300 2.165 8.335 2.335 ;
        RECT 6.045 1.485 6.605 1.575 ;
        RECT 5.725 1.245 6.605 1.485 ;
        RECT 4.905 0.705 5.535 1.035 ;
        RECT 3.725 0.445 3.895 0.695 ;
        RECT 4.565 0.535 4.735 0.695 ;
        RECT 5.725 0.535 5.895 1.245 ;
        RECT 6.775 1.065 6.995 2.135 ;
        RECT 7.165 1.245 7.405 1.965 ;
        RECT 7.575 1.575 7.945 1.905 ;
        RECT 6.065 0.765 6.995 1.065 ;
        RECT 7.575 1.035 7.765 1.575 ;
        RECT 8.165 1.405 8.335 2.165 ;
        RECT 8.565 2.135 8.870 2.635 ;
        RECT 9.220 1.905 9.505 2.455 ;
        RECT 8.555 1.575 9.505 1.905 ;
        RECT 9.690 1.625 9.860 2.635 ;
        RECT 10.670 1.845 10.840 2.635 ;
        RECT 1.535 0.275 1.905 0.445 ;
        RECT 2.125 0.085 2.455 0.445 ;
        RECT 3.070 0.275 3.895 0.445 ;
        RECT 4.115 0.085 4.315 0.525 ;
        RECT 4.565 0.365 4.915 0.535 ;
        RECT 5.135 0.365 5.895 0.535 ;
        RECT 6.225 0.085 6.595 0.585 ;
        RECT 6.775 0.535 6.995 0.765 ;
        RECT 7.165 0.705 7.765 1.035 ;
        RECT 7.985 1.325 8.335 1.405 ;
        RECT 9.320 1.325 9.505 1.575 ;
        RECT 7.985 0.995 9.150 1.325 ;
        RECT 9.320 0.995 10.130 1.325 ;
        RECT 7.985 0.535 8.205 0.995 ;
        RECT 9.320 0.825 9.500 0.995 ;
        RECT 6.775 0.365 7.285 0.535 ;
        RECT 7.565 0.365 8.205 0.535 ;
        RECT 8.450 0.085 8.870 0.615 ;
        RECT 9.140 0.300 9.500 0.825 ;
        RECT 9.690 0.085 9.860 0.695 ;
        RECT 10.670 0.085 10.840 0.565 ;
        RECT 0.000 -0.085 11.040 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 0.665 1.740 0.835 1.910 ;
        RECT 1.155 0.720 1.325 0.890 ;
        RECT 5.665 1.740 5.835 1.910 ;
        RECT 5.155 0.720 5.325 0.890 ;
        RECT 7.225 1.740 7.395 1.910 ;
        RECT 7.225 0.720 7.395 0.890 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
      LAYER met1 ;
        RECT 0.605 1.800 7.455 1.940 ;
        RECT 0.605 1.710 0.895 1.800 ;
        RECT 5.555 1.710 5.895 1.800 ;
        RECT 7.115 1.710 7.455 1.800 ;
        RECT 1.095 0.780 7.455 0.920 ;
        RECT 1.095 0.690 1.385 0.780 ;
        RECT 5.045 0.690 5.385 0.780 ;
        RECT 7.115 0.690 7.455 0.780 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfxtp_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__sdfxtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sdfxtp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.960 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 2.745 1.355 3.150 1.685 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 3.725 1.035 4.095 1.655 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.356400 ;
    PORT
      LAYER li1 ;
        RECT 1.880 0.785 2.215 1.685 ;
        RECT 3.335 0.785 3.505 1.115 ;
        RECT 1.880 0.615 3.505 0.785 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.960 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 6.375 0.785 7.335 1.005 ;
        RECT 9.050 0.785 11.925 1.015 ;
        RECT 0.005 0.725 4.475 0.785 ;
        RECT 5.595 0.725 11.925 0.785 ;
        RECT 0.005 0.105 11.925 0.725 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 12.150 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.960 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.028500 ;
    PORT
      LAYER li1 ;
        RECT 10.030 1.675 10.410 2.395 ;
        RECT 10.980 1.675 11.360 2.395 ;
        RECT 10.030 1.505 11.850 1.675 ;
        RECT 11.550 0.905 11.850 1.505 ;
        RECT 10.030 0.735 11.850 0.905 ;
        RECT 10.030 0.305 10.410 0.735 ;
        RECT 10.980 0.305 11.360 0.735 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 11.960 2.805 ;
        RECT 0.180 1.965 0.350 2.465 ;
        RECT 0.520 2.135 0.900 2.635 ;
        RECT 0.180 1.795 0.895 1.965 ;
        RECT 0.665 0.805 0.895 1.795 ;
        RECT 0.175 0.635 0.895 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.115 0.345 1.345 2.465 ;
        RECT 1.535 2.075 1.810 2.445 ;
        RECT 1.980 2.245 2.360 2.635 ;
        RECT 2.895 2.245 3.890 2.415 ;
        RECT 1.535 1.860 3.525 2.075 ;
        RECT 1.535 0.445 1.705 1.860 ;
        RECT 2.385 1.125 2.555 1.860 ;
        RECT 3.330 1.355 3.525 1.860 ;
        RECT 3.720 1.995 3.890 2.245 ;
        RECT 4.110 2.165 4.280 2.635 ;
        RECT 4.565 2.065 4.800 2.440 ;
        RECT 5.045 2.190 6.265 2.360 ;
        RECT 4.565 1.995 4.735 2.065 ;
        RECT 3.720 1.825 4.735 1.995 ;
        RECT 2.385 0.955 2.715 1.125 ;
        RECT 4.565 0.865 4.735 1.825 ;
        RECT 3.725 0.695 4.735 0.865 ;
        RECT 4.905 1.035 5.195 1.905 ;
        RECT 5.385 1.655 5.875 2.010 ;
        RECT 6.045 1.575 6.265 2.190 ;
        RECT 6.435 1.835 6.605 2.635 ;
        RECT 6.775 2.135 7.075 2.465 ;
        RECT 7.300 2.165 8.335 2.335 ;
        RECT 6.045 1.485 6.605 1.575 ;
        RECT 5.725 1.245 6.605 1.485 ;
        RECT 4.905 0.705 5.535 1.035 ;
        RECT 3.725 0.445 3.895 0.695 ;
        RECT 4.565 0.535 4.735 0.695 ;
        RECT 5.725 0.535 5.895 1.245 ;
        RECT 6.775 1.065 6.995 2.135 ;
        RECT 7.165 1.245 7.405 1.965 ;
        RECT 7.575 1.575 7.945 1.905 ;
        RECT 6.065 0.765 6.995 1.065 ;
        RECT 7.575 1.035 7.765 1.575 ;
        RECT 8.165 1.405 8.335 2.165 ;
        RECT 8.565 2.135 8.870 2.635 ;
        RECT 9.220 1.905 9.505 2.455 ;
        RECT 8.555 1.575 9.505 1.905 ;
        RECT 9.690 1.625 9.860 2.635 ;
        RECT 10.640 1.845 10.810 2.635 ;
        RECT 11.580 1.845 11.750 2.635 ;
        RECT 1.535 0.275 1.905 0.445 ;
        RECT 2.125 0.085 2.455 0.445 ;
        RECT 3.070 0.275 3.895 0.445 ;
        RECT 4.115 0.085 4.315 0.525 ;
        RECT 4.565 0.365 4.915 0.535 ;
        RECT 5.135 0.365 5.895 0.535 ;
        RECT 6.225 0.085 6.595 0.585 ;
        RECT 6.775 0.535 6.995 0.765 ;
        RECT 7.165 0.705 7.765 1.035 ;
        RECT 7.985 1.325 8.335 1.405 ;
        RECT 9.320 1.325 9.505 1.575 ;
        RECT 7.985 0.995 9.150 1.325 ;
        RECT 9.320 1.075 11.380 1.325 ;
        RECT 7.985 0.535 8.205 0.995 ;
        RECT 9.320 0.825 9.500 1.075 ;
        RECT 6.775 0.365 7.285 0.535 ;
        RECT 7.565 0.365 8.205 0.535 ;
        RECT 8.450 0.085 8.870 0.615 ;
        RECT 9.140 0.300 9.500 0.825 ;
        RECT 9.690 0.085 9.860 0.695 ;
        RECT 10.640 0.085 10.810 0.565 ;
        RECT 11.580 0.085 11.750 0.565 ;
        RECT 0.000 -0.085 11.960 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 0.665 1.740 0.835 1.910 ;
        RECT 1.155 0.720 1.325 0.890 ;
        RECT 5.665 1.740 5.835 1.910 ;
        RECT 5.155 0.720 5.325 0.890 ;
        RECT 7.225 1.740 7.395 1.910 ;
        RECT 7.225 0.720 7.395 0.890 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
      LAYER met1 ;
        RECT 0.605 1.800 7.455 1.940 ;
        RECT 0.605 1.710 0.895 1.800 ;
        RECT 5.555 1.710 5.895 1.800 ;
        RECT 7.115 1.710 7.455 1.800 ;
        RECT 1.095 0.780 7.455 0.920 ;
        RECT 1.095 0.690 1.385 0.780 ;
        RECT 5.045 0.690 5.385 0.780 ;
        RECT 7.115 0.690 7.455 0.780 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfxtp_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__sdlclkp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sdlclkp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.356400 ;
    PORT
      LAYER met1 ;
        RECT 4.745 1.260 5.035 1.305 ;
        RECT 5.940 1.260 6.230 1.305 ;
        RECT 4.745 1.120 6.230 1.260 ;
        RECT 4.745 1.075 5.035 1.120 ;
        RECT 5.940 1.075 6.230 1.120 ;
    END
  END CLK
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.855 0.955 1.235 1.955 ;
    END
  END GATE
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.955 0.330 1.665 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.720 0.785 3.715 1.015 ;
        RECT 6.330 0.785 7.325 1.015 ;
        RECT 0.005 0.105 7.325 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.480250 ;
    PORT
      LAYER li1 ;
        RECT 6.985 0.255 7.235 2.465 ;
    END
  END GCLK
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.360 2.805 ;
        RECT 0.085 1.835 0.345 2.635 ;
        RECT 0.515 2.125 1.280 2.465 ;
        RECT 1.610 2.125 2.300 2.465 ;
        RECT 0.515 0.785 0.685 2.125 ;
        RECT 1.465 1.205 1.960 1.955 ;
        RECT 2.130 1.375 2.300 2.125 ;
        RECT 2.520 2.075 3.105 2.635 ;
        RECT 3.325 2.085 3.545 2.465 ;
        RECT 3.885 2.255 5.735 2.635 ;
        RECT 5.955 2.085 6.125 2.465 ;
        RECT 6.385 2.255 6.715 2.635 ;
        RECT 3.325 1.915 5.735 2.085 ;
        RECT 3.325 1.905 3.545 1.915 ;
        RECT 2.470 1.635 3.545 1.905 ;
        RECT 2.470 1.575 2.665 1.635 ;
        RECT 2.130 1.205 3.205 1.375 ;
        RECT 0.085 0.615 1.295 0.785 ;
        RECT 1.465 0.705 1.800 1.205 ;
        RECT 1.970 0.705 2.305 1.035 ;
        RECT 2.475 0.995 3.205 1.205 ;
        RECT 0.085 0.255 0.345 0.615 ;
        RECT 0.515 0.085 0.895 0.445 ;
        RECT 1.115 0.255 1.295 0.615 ;
        RECT 2.475 0.535 2.645 0.995 ;
        RECT 1.465 0.255 2.645 0.535 ;
        RECT 2.910 0.085 3.080 0.825 ;
        RECT 3.375 0.255 3.545 1.635 ;
        RECT 3.735 1.575 4.145 1.745 ;
        RECT 3.735 0.935 3.905 1.575 ;
        RECT 4.365 1.495 5.215 1.745 ;
        RECT 4.365 1.275 4.550 1.495 ;
        RECT 4.075 1.105 4.550 1.275 ;
        RECT 3.735 0.255 4.065 0.935 ;
        RECT 4.380 0.785 4.550 1.105 ;
        RECT 4.745 0.995 5.060 1.325 ;
        RECT 5.385 0.995 5.735 1.915 ;
        RECT 5.955 1.495 6.815 2.085 ;
        RECT 5.955 0.995 6.395 1.325 ;
        RECT 6.645 0.785 6.815 1.495 ;
        RECT 4.380 0.615 5.215 0.785 ;
        RECT 4.285 0.085 4.615 0.445 ;
        RECT 4.965 0.255 5.215 0.615 ;
        RECT 5.535 0.615 6.815 0.785 ;
        RECT 5.535 0.255 5.705 0.615 ;
        RECT 6.325 0.085 6.685 0.445 ;
        RECT 0.000 -0.085 7.360 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 1.625 1.445 1.795 1.615 ;
        RECT 2.135 0.765 2.305 0.935 ;
        RECT 4.365 1.445 4.535 1.615 ;
        RECT 3.800 0.765 3.970 0.935 ;
        RECT 4.805 1.105 4.975 1.275 ;
        RECT 6.000 1.105 6.170 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
      LAYER met1 ;
        RECT 1.565 1.600 1.855 1.645 ;
        RECT 4.305 1.600 4.595 1.645 ;
        RECT 1.565 1.460 4.595 1.600 ;
        RECT 1.565 1.415 1.855 1.460 ;
        RECT 4.305 1.415 4.595 1.460 ;
        RECT 2.075 0.920 2.365 0.965 ;
        RECT 3.740 0.920 4.030 0.965 ;
        RECT 2.075 0.780 4.030 0.920 ;
        RECT 2.075 0.735 2.365 0.780 ;
        RECT 3.740 0.735 4.030 0.780 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdlclkp_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__sdlclkp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sdlclkp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.820 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.356400 ;
    PORT
      LAYER met1 ;
        RECT 4.950 1.260 5.240 1.305 ;
        RECT 5.940 1.260 6.230 1.305 ;
        RECT 4.950 1.120 6.230 1.260 ;
        RECT 4.950 1.075 5.240 1.120 ;
        RECT 5.940 1.075 6.230 1.120 ;
    END
  END CLK
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.890 0.955 1.295 1.955 ;
    END
  END GATE
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.955 0.330 1.665 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.820 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.720 0.785 3.715 1.015 ;
        RECT 6.230 0.785 7.730 1.015 ;
        RECT 0.005 0.105 7.730 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.010 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.820 2.960 ;
    END
  END VPWR
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.498000 ;
    PORT
      LAYER li1 ;
        RECT 6.970 1.655 7.220 2.465 ;
        RECT 6.970 1.485 7.675 1.655 ;
        RECT 7.490 0.885 7.675 1.485 ;
        RECT 6.970 0.715 7.675 0.885 ;
        RECT 6.970 0.445 7.170 0.715 ;
        RECT 6.840 0.255 7.170 0.445 ;
    END
  END GCLK
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.820 2.805 ;
        RECT 0.085 1.835 0.345 2.635 ;
        RECT 0.515 2.125 1.280 2.465 ;
        RECT 1.610 2.125 2.300 2.465 ;
        RECT 0.515 0.785 0.720 2.125 ;
        RECT 1.465 1.205 1.960 1.955 ;
        RECT 2.130 1.375 2.300 2.125 ;
        RECT 2.520 2.075 3.105 2.635 ;
        RECT 3.325 2.085 3.545 2.465 ;
        RECT 3.885 2.255 5.755 2.635 ;
        RECT 5.975 2.085 6.145 2.465 ;
        RECT 6.395 2.255 6.725 2.635 ;
        RECT 3.325 1.915 5.755 2.085 ;
        RECT 3.325 1.905 3.545 1.915 ;
        RECT 2.470 1.635 3.545 1.905 ;
        RECT 2.470 1.575 2.665 1.635 ;
        RECT 2.130 1.205 3.205 1.375 ;
        RECT 0.085 0.615 1.295 0.785 ;
        RECT 1.465 0.705 1.800 1.205 ;
        RECT 1.970 0.705 2.305 1.035 ;
        RECT 2.475 0.995 3.205 1.205 ;
        RECT 0.085 0.255 0.345 0.615 ;
        RECT 0.515 0.085 0.895 0.445 ;
        RECT 1.115 0.255 1.295 0.615 ;
        RECT 2.475 0.535 2.645 0.995 ;
        RECT 1.465 0.255 2.645 0.535 ;
        RECT 2.910 0.085 3.080 0.825 ;
        RECT 3.375 0.255 3.545 1.635 ;
        RECT 3.735 1.575 4.145 1.745 ;
        RECT 3.735 0.935 3.905 1.575 ;
        RECT 4.365 1.495 5.215 1.745 ;
        RECT 4.365 1.275 4.670 1.495 ;
        RECT 4.075 1.105 4.670 1.275 ;
        RECT 3.735 0.765 4.160 0.935 ;
        RECT 4.380 0.785 4.670 1.105 ;
        RECT 4.965 0.995 5.185 1.325 ;
        RECT 5.405 0.995 5.755 1.915 ;
        RECT 5.975 1.495 6.750 2.085 ;
        RECT 7.440 1.825 7.690 2.635 ;
        RECT 5.975 0.995 6.405 1.325 ;
        RECT 6.580 1.315 6.750 1.495 ;
        RECT 6.580 1.055 7.270 1.315 ;
        RECT 6.580 0.785 6.750 1.055 ;
        RECT 3.735 0.255 4.065 0.765 ;
        RECT 4.380 0.615 5.085 0.785 ;
        RECT 4.285 0.085 4.615 0.445 ;
        RECT 4.835 0.255 5.085 0.615 ;
        RECT 5.505 0.615 6.750 0.785 ;
        RECT 5.505 0.255 5.675 0.615 ;
        RECT 6.335 0.085 6.670 0.445 ;
        RECT 7.390 0.085 7.560 0.545 ;
        RECT 0.000 -0.085 7.820 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 1.625 1.445 1.795 1.615 ;
        RECT 2.135 0.765 2.305 0.935 ;
        RECT 4.500 1.445 4.670 1.615 ;
        RECT 3.990 0.765 4.160 0.935 ;
        RECT 5.010 1.105 5.180 1.275 ;
        RECT 6.000 1.105 6.170 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
      LAYER met1 ;
        RECT 1.565 1.600 1.855 1.645 ;
        RECT 4.440 1.600 4.730 1.645 ;
        RECT 1.565 1.460 4.730 1.600 ;
        RECT 1.565 1.415 1.855 1.460 ;
        RECT 4.440 1.415 4.730 1.460 ;
        RECT 2.075 0.920 2.365 0.965 ;
        RECT 3.930 0.920 4.220 0.965 ;
        RECT 2.075 0.780 4.220 0.920 ;
        RECT 2.075 0.735 2.365 0.780 ;
        RECT 3.930 0.735 4.220 0.780 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdlclkp_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__sdlclkp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sdlclkp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.200 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.455700 ;
    PORT
      LAYER met1 ;
        RECT 5.055 1.260 5.345 1.305 ;
        RECT 6.100 1.260 6.390 1.305 ;
        RECT 5.055 1.120 6.390 1.260 ;
        RECT 5.055 1.075 5.345 1.120 ;
        RECT 6.100 1.075 6.390 1.120 ;
    END
  END CLK
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.905 1.445 1.340 1.955 ;
        RECT 0.905 0.955 1.295 1.445 ;
    END
  END GATE
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.955 0.345 1.665 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.200 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.780 0.785 3.875 1.015 ;
        RECT 5.495 0.785 9.125 1.015 ;
        RECT 0.005 0.105 9.125 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.390 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.200 2.960 ;
    END
  END VPWR
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.251250 ;
    PORT
      LAYER li1 ;
        RECT 7.130 1.655 7.380 2.465 ;
        RECT 7.130 1.485 7.820 1.655 ;
        RECT 7.650 1.315 7.820 1.485 ;
        RECT 8.205 1.315 8.595 2.465 ;
        RECT 7.650 1.055 9.055 1.315 ;
        RECT 7.650 0.885 7.820 1.055 ;
        RECT 7.130 0.715 7.820 0.885 ;
        RECT 7.130 0.445 7.380 0.715 ;
        RECT 7.000 0.255 7.380 0.445 ;
        RECT 8.205 0.255 8.595 1.055 ;
    END
  END GCLK
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.200 2.805 ;
        RECT 0.085 1.835 0.345 2.635 ;
        RECT 0.515 2.125 1.360 2.465 ;
        RECT 1.530 2.125 2.405 2.465 ;
        RECT 0.515 0.785 0.735 2.125 ;
        RECT 1.510 1.325 2.015 1.955 ;
        RECT 1.465 1.205 2.015 1.325 ;
        RECT 2.235 1.375 2.405 2.125 ;
        RECT 2.575 2.075 3.265 2.635 ;
        RECT 3.485 2.085 3.705 2.465 ;
        RECT 3.895 2.255 5.915 2.635 ;
        RECT 6.135 2.085 6.305 2.465 ;
        RECT 6.555 2.255 6.885 2.635 ;
        RECT 3.485 1.915 5.915 2.085 ;
        RECT 3.485 1.905 3.705 1.915 ;
        RECT 2.575 1.635 3.705 1.905 ;
        RECT 2.575 1.575 2.795 1.635 ;
        RECT 2.235 1.205 3.265 1.375 ;
        RECT 0.085 0.615 1.295 0.785 ;
        RECT 1.465 0.705 1.855 1.205 ;
        RECT 2.025 0.705 2.360 1.035 ;
        RECT 2.530 0.995 3.265 1.205 ;
        RECT 0.085 0.255 0.345 0.615 ;
        RECT 0.515 0.085 0.895 0.445 ;
        RECT 1.115 0.255 1.295 0.615 ;
        RECT 2.530 0.535 2.700 0.995 ;
        RECT 1.465 0.255 2.700 0.535 ;
        RECT 2.920 0.085 3.265 0.825 ;
        RECT 3.485 0.255 3.705 1.635 ;
        RECT 3.895 1.575 4.305 1.745 ;
        RECT 3.895 0.935 4.065 1.575 ;
        RECT 4.525 1.495 5.375 1.745 ;
        RECT 4.525 1.275 4.830 1.495 ;
        RECT 4.235 1.105 4.830 1.275 ;
        RECT 3.895 0.765 4.320 0.935 ;
        RECT 4.540 0.785 4.830 1.105 ;
        RECT 5.055 0.995 5.345 1.325 ;
        RECT 5.565 0.995 5.915 1.915 ;
        RECT 6.135 1.495 6.910 2.085 ;
        RECT 7.600 1.825 7.850 2.635 ;
        RECT 6.135 0.995 6.565 1.325 ;
        RECT 6.740 1.315 6.910 1.495 ;
        RECT 8.765 1.485 9.035 2.635 ;
        RECT 6.740 1.055 7.430 1.315 ;
        RECT 6.740 0.785 6.910 1.055 ;
        RECT 3.895 0.255 4.225 0.765 ;
        RECT 4.540 0.615 5.245 0.785 ;
        RECT 4.395 0.085 4.775 0.445 ;
        RECT 4.995 0.255 5.245 0.615 ;
        RECT 5.415 0.615 6.910 0.785 ;
        RECT 5.415 0.255 5.835 0.615 ;
        RECT 6.005 0.085 6.830 0.445 ;
        RECT 7.600 0.085 7.850 0.545 ;
        RECT 8.765 0.085 9.035 0.885 ;
        RECT 0.000 -0.085 9.200 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 1.680 1.445 1.850 1.615 ;
        RECT 2.190 0.765 2.360 0.935 ;
        RECT 4.660 1.445 4.830 1.615 ;
        RECT 4.150 0.765 4.320 0.935 ;
        RECT 5.115 1.105 5.285 1.275 ;
        RECT 6.160 1.105 6.330 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
      LAYER met1 ;
        RECT 1.620 1.600 1.910 1.645 ;
        RECT 4.600 1.600 4.890 1.645 ;
        RECT 1.620 1.460 4.890 1.600 ;
        RECT 1.620 1.415 1.910 1.460 ;
        RECT 4.600 1.415 4.890 1.460 ;
        RECT 2.130 0.920 2.420 0.965 ;
        RECT 4.090 0.920 4.380 0.965 ;
        RECT 2.130 0.780 4.380 0.920 ;
        RECT 2.130 0.735 2.420 0.780 ;
        RECT 4.090 0.735 4.380 0.780 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdlclkp_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__sedfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sedfxbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.180 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 1.795 0.765 2.155 1.720 ;
    END
  END D
  PIN DE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.356400 ;
    PORT
      LAYER li1 ;
        RECT 2.325 1.185 2.525 1.370 ;
        RECT 2.325 0.765 2.765 1.185 ;
    END
  END DE
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 6.445 1.105 6.950 1.665 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.356400 ;
    PORT
      LAYER li1 ;
        RECT 5.605 1.105 5.885 1.615 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 15.180 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 5.805 0.785 7.920 1.145 ;
        RECT 9.335 0.785 10.305 1.005 ;
        RECT 12.450 0.785 15.085 1.015 ;
        RECT 0.005 0.465 15.085 0.785 ;
        RECT 0.005 0.105 5.365 0.465 ;
        RECT 7.220 0.105 15.085 0.465 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.435 15.370 2.910 ;
        RECT -0.190 1.305 5.285 1.435 ;
        RECT 7.985 1.305 15.370 1.435 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 15.180 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.513250 ;
    PORT
      LAYER li1 ;
        RECT 14.655 0.255 15.070 2.420 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 12.960 0.255 13.315 2.465 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 15.180 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.895 2.635 ;
        RECT 0.175 1.795 0.895 1.965 ;
        RECT 0.665 0.805 0.895 1.795 ;
        RECT 0.175 0.635 0.895 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.115 0.345 1.285 2.465 ;
        RECT 1.455 1.890 1.885 2.465 ;
        RECT 2.385 1.890 2.765 2.635 ;
        RECT 1.455 0.515 1.625 1.890 ;
        RECT 2.955 1.720 3.285 2.425 ;
        RECT 3.515 1.825 3.710 2.635 ;
        RECT 4.425 2.020 4.805 2.465 ;
        RECT 5.035 2.210 5.365 2.465 ;
        RECT 4.425 1.820 4.865 2.020 ;
        RECT 2.695 1.355 3.285 1.720 ;
        RECT 2.980 1.175 3.285 1.355 ;
        RECT 4.105 1.320 4.525 1.650 ;
        RECT 2.980 0.845 3.885 1.175 ;
        RECT 1.455 0.255 1.885 0.515 ;
        RECT 2.385 0.085 2.765 0.515 ;
        RECT 2.980 0.255 3.205 0.845 ;
        RECT 4.105 0.685 4.275 1.320 ;
        RECT 4.695 1.150 4.865 1.820 ;
        RECT 4.445 0.980 4.865 1.150 ;
        RECT 5.085 1.785 5.365 2.210 ;
        RECT 5.790 2.005 6.130 2.465 ;
        RECT 6.350 2.175 6.695 2.635 ;
        RECT 7.460 2.150 7.790 2.465 ;
        RECT 8.000 2.175 9.190 2.375 ;
        RECT 5.790 1.835 7.370 2.005 ;
        RECT 3.385 0.085 3.765 0.610 ;
        RECT 4.445 0.255 4.765 0.980 ;
        RECT 5.085 0.825 5.255 1.785 ;
        RECT 6.055 0.935 6.225 1.835 ;
        RECT 7.120 1.355 7.370 1.835 ;
        RECT 7.540 1.865 7.790 2.150 ;
        RECT 7.540 1.185 7.710 1.865 ;
        RECT 4.995 0.645 5.255 0.825 ;
        RECT 4.995 0.255 5.195 0.645 ;
        RECT 5.895 0.515 6.225 0.935 ;
        RECT 5.365 0.255 6.225 0.515 ;
        RECT 6.445 0.085 6.695 0.905 ;
        RECT 7.300 0.565 7.710 1.185 ;
        RECT 7.880 1.125 8.115 1.720 ;
        RECT 8.285 1.655 8.800 2.005 ;
        RECT 8.285 0.955 8.455 1.655 ;
        RECT 8.970 1.575 9.190 2.175 ;
        RECT 9.360 1.835 9.595 2.635 ;
        RECT 8.970 1.485 9.595 1.575 ;
        RECT 7.900 0.735 8.455 0.955 ;
        RECT 8.695 1.315 9.595 1.485 ;
        RECT 8.695 0.565 8.865 1.315 ;
        RECT 9.425 1.245 9.595 1.315 ;
        RECT 9.765 1.375 10.145 2.465 ;
        RECT 10.355 2.105 10.645 2.635 ;
        RECT 11.260 2.165 12.375 2.355 ;
        RECT 9.055 1.065 9.305 1.095 ;
        RECT 9.765 1.065 10.730 1.375 ;
        RECT 11.125 1.245 11.365 1.965 ;
        RECT 9.055 1.045 10.730 1.065 ;
        RECT 9.055 0.765 10.220 1.045 ;
        RECT 11.535 1.035 11.905 1.995 ;
        RECT 7.300 0.255 7.920 0.565 ;
        RECT 8.140 0.255 8.865 0.565 ;
        RECT 9.180 0.085 9.575 0.560 ;
        RECT 9.765 0.255 10.220 0.765 ;
        RECT 11.375 0.705 11.905 1.035 ;
        RECT 10.450 0.085 10.725 0.615 ;
        RECT 12.125 0.535 12.375 2.165 ;
        RECT 12.595 1.495 12.765 2.635 ;
        RECT 13.605 1.220 13.945 2.465 ;
        RECT 14.165 1.465 14.400 2.635 ;
        RECT 11.410 0.330 12.375 0.535 ;
        RECT 12.545 0.085 12.790 0.900 ;
        RECT 13.485 0.890 13.945 1.220 ;
        RECT 14.115 1.070 14.445 1.295 ;
        RECT 13.605 0.255 13.945 0.890 ;
        RECT 14.165 0.085 14.400 0.900 ;
        RECT 0.000 -0.085 15.180 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 14.405 2.635 14.575 2.805 ;
        RECT 14.865 2.635 15.035 2.805 ;
        RECT 0.685 1.785 0.855 1.955 ;
        RECT 1.115 1.445 1.285 1.615 ;
        RECT 1.455 0.425 1.625 0.595 ;
        RECT 4.105 0.765 4.275 0.935 ;
        RECT 8.345 1.785 8.515 1.955 ;
        RECT 4.535 0.425 4.705 0.595 ;
        RECT 5.015 0.425 5.185 0.595 ;
        RECT 7.910 1.445 8.080 1.615 ;
        RECT 7.315 0.425 7.485 0.595 ;
        RECT 11.160 1.785 11.330 1.955 ;
        RECT 11.630 1.445 11.800 1.615 ;
        RECT 12.165 1.105 12.335 1.275 ;
        RECT 14.195 1.105 14.365 1.275 ;
        RECT 13.700 0.765 13.870 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
        RECT 14.405 -0.085 14.575 0.085 ;
        RECT 14.865 -0.085 15.035 0.085 ;
      LAYER met1 ;
        RECT 0.625 1.940 0.915 1.985 ;
        RECT 8.285 1.940 8.625 1.985 ;
        RECT 11.075 1.940 11.415 1.985 ;
        RECT 0.625 1.800 11.415 1.940 ;
        RECT 0.625 1.755 0.915 1.800 ;
        RECT 8.285 1.755 8.625 1.800 ;
        RECT 11.075 1.755 11.415 1.800 ;
        RECT 1.005 1.600 1.345 1.645 ;
        RECT 7.825 1.600 8.165 1.645 ;
        RECT 11.545 1.600 11.885 1.645 ;
        RECT 1.005 1.460 11.885 1.600 ;
        RECT 1.005 1.415 1.345 1.460 ;
        RECT 7.825 1.415 8.165 1.460 ;
        RECT 11.545 1.415 11.885 1.460 ;
        RECT 12.105 1.260 12.395 1.305 ;
        RECT 14.135 1.260 14.425 1.305 ;
        RECT 12.105 1.120 14.425 1.260 ;
        RECT 12.105 1.075 12.395 1.120 ;
        RECT 14.135 1.075 14.425 1.120 ;
        RECT 4.045 0.920 4.335 0.965 ;
        RECT 13.640 0.920 13.930 0.965 ;
        RECT 4.045 0.780 13.930 0.920 ;
        RECT 4.045 0.735 4.335 0.780 ;
        RECT 13.640 0.735 13.930 0.780 ;
        RECT 1.395 0.580 1.685 0.625 ;
        RECT 4.425 0.580 4.765 0.625 ;
        RECT 1.395 0.395 4.765 0.580 ;
        RECT 4.905 0.580 5.245 0.625 ;
        RECT 7.205 0.580 7.545 0.625 ;
        RECT 4.905 0.395 7.545 0.580 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sedfxbp_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__sedfxbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sedfxbp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.560 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 1.795 0.765 2.155 1.720 ;
    END
  END D
  PIN DE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.356400 ;
    PORT
      LAYER li1 ;
        RECT 2.325 1.185 2.525 1.370 ;
        RECT 2.325 0.765 2.765 1.185 ;
    END
  END DE
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.178200 ;
    PORT
      LAYER li1 ;
        RECT 6.445 1.105 6.950 1.665 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.356400 ;
    PORT
      LAYER li1 ;
        RECT 5.605 1.105 5.885 1.615 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 16.560 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 5.805 0.785 7.920 1.145 ;
        RECT 9.335 0.785 10.305 1.005 ;
        RECT 12.540 0.785 16.280 1.015 ;
        RECT 0.005 0.465 16.280 0.785 ;
        RECT 0.005 0.105 5.365 0.465 ;
        RECT 7.220 0.105 16.280 0.465 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.435 16.750 2.910 ;
        RECT -0.190 1.305 5.285 1.435 ;
        RECT 7.985 1.305 16.750 1.435 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 16.560 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.530500 ;
    PORT
      LAYER li1 ;
        RECT 15.320 0.255 15.700 2.420 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.498000 ;
    PORT
      LAYER li1 ;
        RECT 12.935 1.300 13.315 2.465 ;
        RECT 12.935 1.065 13.430 1.300 ;
        RECT 13.100 0.255 13.430 1.065 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 16.560 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.895 2.635 ;
        RECT 0.175 1.795 0.895 1.965 ;
        RECT 0.665 0.805 0.895 1.795 ;
        RECT 0.175 0.635 0.895 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.895 0.465 ;
        RECT 1.115 0.345 1.285 2.465 ;
        RECT 1.455 1.890 1.885 2.465 ;
        RECT 2.385 1.890 2.765 2.635 ;
        RECT 1.455 0.515 1.625 1.890 ;
        RECT 2.955 1.720 3.285 2.425 ;
        RECT 3.515 1.825 3.710 2.635 ;
        RECT 4.425 2.020 4.805 2.465 ;
        RECT 5.035 2.210 5.365 2.465 ;
        RECT 4.425 1.820 4.865 2.020 ;
        RECT 2.695 1.355 3.285 1.720 ;
        RECT 2.980 1.175 3.285 1.355 ;
        RECT 4.105 1.320 4.525 1.650 ;
        RECT 2.980 0.845 3.885 1.175 ;
        RECT 1.455 0.255 1.885 0.515 ;
        RECT 2.385 0.085 2.765 0.515 ;
        RECT 2.980 0.255 3.205 0.845 ;
        RECT 4.105 0.685 4.275 1.320 ;
        RECT 4.695 1.150 4.865 1.820 ;
        RECT 4.445 0.980 4.865 1.150 ;
        RECT 5.085 1.785 5.365 2.210 ;
        RECT 5.790 2.005 6.130 2.465 ;
        RECT 6.350 2.175 6.695 2.635 ;
        RECT 7.460 2.150 7.790 2.465 ;
        RECT 8.000 2.175 9.190 2.375 ;
        RECT 5.790 1.835 7.370 2.005 ;
        RECT 3.385 0.085 3.765 0.610 ;
        RECT 4.445 0.255 4.765 0.980 ;
        RECT 5.085 0.825 5.255 1.785 ;
        RECT 6.055 0.935 6.225 1.835 ;
        RECT 7.120 1.355 7.370 1.835 ;
        RECT 7.540 1.865 7.790 2.150 ;
        RECT 7.540 1.185 7.710 1.865 ;
        RECT 4.995 0.645 5.255 0.825 ;
        RECT 4.995 0.255 5.195 0.645 ;
        RECT 5.895 0.515 6.225 0.935 ;
        RECT 5.365 0.255 6.225 0.515 ;
        RECT 6.445 0.085 6.695 0.905 ;
        RECT 7.300 0.565 7.710 1.185 ;
        RECT 7.880 1.125 8.115 1.720 ;
        RECT 8.285 1.655 8.800 2.005 ;
        RECT 8.285 0.955 8.455 1.655 ;
        RECT 8.970 1.575 9.190 2.175 ;
        RECT 9.360 1.835 9.595 2.635 ;
        RECT 8.970 1.485 9.595 1.575 ;
        RECT 7.900 0.735 8.455 0.955 ;
        RECT 8.695 1.315 9.595 1.485 ;
        RECT 8.695 0.565 8.865 1.315 ;
        RECT 9.425 1.245 9.595 1.315 ;
        RECT 9.765 1.375 10.145 2.465 ;
        RECT 10.355 2.105 10.645 2.635 ;
        RECT 11.260 2.165 12.375 2.355 ;
        RECT 9.055 1.065 9.305 1.095 ;
        RECT 9.765 1.065 10.730 1.375 ;
        RECT 11.125 1.245 11.365 1.965 ;
        RECT 9.055 1.045 10.730 1.065 ;
        RECT 9.055 0.765 10.220 1.045 ;
        RECT 11.535 1.035 11.905 1.995 ;
        RECT 7.300 0.255 7.920 0.565 ;
        RECT 8.140 0.255 8.865 0.565 ;
        RECT 9.180 0.085 9.575 0.560 ;
        RECT 9.765 0.255 10.220 0.765 ;
        RECT 11.390 0.705 11.905 1.035 ;
        RECT 10.450 0.085 10.725 0.615 ;
        RECT 12.125 0.535 12.375 2.165 ;
        RECT 12.595 1.495 12.765 2.635 ;
        RECT 13.535 1.465 13.785 2.635 ;
        RECT 13.955 1.575 14.185 2.010 ;
        RECT 14.355 1.220 14.695 2.465 ;
        RECT 14.915 1.465 15.150 2.635 ;
        RECT 15.920 1.465 16.180 2.635 ;
        RECT 11.410 0.330 12.375 0.535 ;
        RECT 12.630 0.085 12.880 0.900 ;
        RECT 13.650 0.085 13.900 0.900 ;
        RECT 14.070 0.890 14.695 1.220 ;
        RECT 14.355 0.255 14.695 0.890 ;
        RECT 14.915 0.085 15.150 0.900 ;
        RECT 15.920 0.085 16.180 0.900 ;
        RECT 0.000 -0.085 16.560 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 14.405 2.635 14.575 2.805 ;
        RECT 14.865 2.635 15.035 2.805 ;
        RECT 15.325 2.635 15.495 2.805 ;
        RECT 15.785 2.635 15.955 2.805 ;
        RECT 16.245 2.635 16.415 2.805 ;
        RECT 0.685 1.785 0.855 1.955 ;
        RECT 1.115 1.445 1.285 1.615 ;
        RECT 1.455 0.425 1.625 0.595 ;
        RECT 4.105 0.765 4.275 0.935 ;
        RECT 8.345 1.785 8.515 1.955 ;
        RECT 4.535 0.425 4.705 0.595 ;
        RECT 5.015 0.425 5.185 0.595 ;
        RECT 7.910 1.445 8.080 1.615 ;
        RECT 7.315 0.425 7.485 0.595 ;
        RECT 11.160 1.785 11.330 1.955 ;
        RECT 11.630 1.445 11.800 1.615 ;
        RECT 12.165 1.785 12.335 1.955 ;
        RECT 13.985 1.785 14.155 1.955 ;
        RECT 14.445 0.765 14.615 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
        RECT 14.405 -0.085 14.575 0.085 ;
        RECT 14.865 -0.085 15.035 0.085 ;
        RECT 15.325 -0.085 15.495 0.085 ;
        RECT 15.785 -0.085 15.955 0.085 ;
        RECT 16.245 -0.085 16.415 0.085 ;
      LAYER met1 ;
        RECT 0.625 1.940 0.915 1.985 ;
        RECT 8.285 1.940 8.625 1.985 ;
        RECT 11.075 1.940 11.415 1.985 ;
        RECT 0.625 1.800 11.415 1.940 ;
        RECT 0.625 1.755 0.915 1.800 ;
        RECT 8.285 1.755 8.625 1.800 ;
        RECT 11.075 1.755 11.415 1.800 ;
        RECT 12.105 1.940 12.395 1.985 ;
        RECT 13.925 1.940 14.215 1.985 ;
        RECT 12.105 1.800 14.215 1.940 ;
        RECT 12.105 1.755 12.395 1.800 ;
        RECT 13.925 1.755 14.215 1.800 ;
        RECT 1.005 1.600 1.345 1.645 ;
        RECT 7.825 1.600 8.165 1.645 ;
        RECT 11.545 1.600 11.885 1.645 ;
        RECT 1.005 1.460 11.885 1.600 ;
        RECT 1.005 1.415 1.345 1.460 ;
        RECT 7.825 1.415 8.165 1.460 ;
        RECT 11.545 1.415 11.885 1.460 ;
        RECT 4.045 0.920 4.335 0.965 ;
        RECT 14.385 0.920 14.675 0.965 ;
        RECT 4.045 0.780 14.675 0.920 ;
        RECT 4.045 0.735 4.335 0.780 ;
        RECT 14.385 0.735 14.675 0.780 ;
        RECT 1.395 0.580 1.685 0.625 ;
        RECT 4.425 0.580 4.765 0.625 ;
        RECT 1.395 0.395 4.765 0.580 ;
        RECT 4.905 0.580 5.245 0.625 ;
        RECT 7.205 0.580 7.545 0.625 ;
        RECT 4.905 0.395 7.545 0.580 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sedfxbp_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__tap_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hdll__tap_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.460 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 0.460 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.015 0.190 0.445 0.975 ;
      LAYER li1 ;
        RECT 0.085 0.265 0.375 0.810 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 0.650 2.910 ;
      LAYER li1 ;
        RECT 0.085 1.470 0.375 2.455 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 0.460 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 0.460 2.805 ;
        RECT 0.000 -0.085 0.460 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__tap_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__tapvgnd2_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hdll__tapvgnd2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.460 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.015 0.190 0.445 0.975 ;
      LAYER met1 ;
        RECT 0.000 -0.240 0.460 0.240 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 0.650 2.910 ;
      LAYER met1 ;
        RECT 0.085 1.755 0.375 1.985 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 0.460 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 0.460 2.805 ;
        RECT 0.085 1.470 0.375 2.455 ;
        RECT 0.085 0.085 0.375 0.810 ;
        RECT 0.000 -0.085 0.460 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.145 1.785 0.315 1.955 ;
        RECT 0.145 -0.085 0.315 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__tapvgnd2_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__tapvgnd_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hdll__tapvgnd_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.460 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.015 0.190 0.445 0.975 ;
      LAYER met1 ;
        RECT 0.000 -0.240 0.460 0.240 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 0.650 2.910 ;
      LAYER met1 ;
        RECT 0.085 2.095 0.375 2.325 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 0.460 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 0.460 2.805 ;
        RECT 0.085 1.470 0.375 2.455 ;
        RECT 0.085 0.085 0.375 0.810 ;
        RECT 0.000 -0.085 0.460 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.145 2.125 0.315 2.295 ;
        RECT 0.145 -0.085 0.315 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__tapvgnd_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__tapvpwrvgnd_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hdll__tapvpwrvgnd_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.460 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.015 0.190 0.445 0.975 ;
      LAYER met1 ;
        RECT 0.000 -0.240 0.460 0.240 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 0.650 2.910 ;
      LAYER met1 ;
        RECT 0.000 2.480 0.460 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 0.460 2.805 ;
        RECT 0.085 1.470 0.375 2.635 ;
        RECT 0.085 0.085 0.375 0.810 ;
        RECT 0.000 -0.085 0.460 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__tapvpwrvgnd_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__xnor2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__xnor2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.980 1.075 1.775 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.445 2.165 1.615 ;
        RECT 0.425 0.995 0.810 1.445 ;
        RECT 1.945 1.245 2.165 1.445 ;
        RECT 1.945 1.075 2.645 1.245 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.105 0.105 3.515 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.545000 ;
    PORT
      LAYER li1 ;
        RECT 2.515 2.125 2.895 2.295 ;
        RECT 2.725 1.955 2.895 2.125 ;
        RECT 2.725 1.755 3.595 1.955 ;
        RECT 3.355 0.825 3.595 1.755 ;
        RECT 3.175 0.345 3.595 0.825 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.085 2.125 0.385 2.635 ;
        RECT 0.555 1.955 0.935 2.465 ;
        RECT 1.155 2.125 1.835 2.635 ;
        RECT 3.115 2.125 3.415 2.635 ;
        RECT 0.085 1.785 2.555 1.955 ;
        RECT 0.085 0.825 0.255 1.785 ;
        RECT 2.335 1.585 2.555 1.785 ;
        RECT 2.335 1.415 3.095 1.585 ;
        RECT 2.875 0.995 3.095 1.415 ;
        RECT 0.085 0.280 0.550 0.825 ;
        RECT 1.155 0.085 1.325 0.905 ;
        RECT 1.495 0.655 2.895 0.825 ;
        RECT 1.495 0.255 1.875 0.655 ;
        RECT 2.095 0.085 2.495 0.475 ;
        RECT 2.665 0.255 2.895 0.655 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xnor2_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__xnor2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__xnor2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 1.355 1.075 2.905 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.840 1.445 3.350 1.615 ;
        RECT 0.840 1.285 1.010 1.445 ;
        RECT 0.485 1.075 1.010 1.285 ;
        RECT 3.180 1.285 3.350 1.445 ;
        RECT 3.180 1.075 4.305 1.285 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 6.345 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.953000 ;
    PORT
      LAYER li1 ;
        RECT 4.075 1.965 4.285 2.125 ;
        RECT 5.495 1.965 5.745 2.125 ;
        RECT 4.075 1.795 5.745 1.965 ;
        RECT 5.495 1.625 5.745 1.795 ;
        RECT 5.495 1.415 6.340 1.625 ;
        RECT 5.950 0.475 6.340 1.415 ;
        RECT 4.985 0.305 6.340 0.475 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.085 1.965 0.400 2.465 ;
        RECT 0.620 2.135 0.870 2.635 ;
        RECT 1.090 1.965 1.340 2.465 ;
        RECT 1.560 2.135 1.810 2.635 ;
        RECT 2.030 1.965 2.280 2.465 ;
        RECT 2.590 2.125 2.840 2.465 ;
        RECT 3.060 2.135 3.310 2.635 ;
        RECT 3.530 2.295 4.755 2.465 ;
        RECT 3.530 2.125 3.855 2.295 ;
        RECT 4.505 2.135 4.755 2.295 ;
        RECT 5.025 2.135 5.275 2.635 ;
        RECT 0.085 1.955 2.280 1.965 ;
        RECT 0.085 1.785 3.780 1.955 ;
        RECT 5.965 1.795 6.340 2.635 ;
        RECT 0.085 0.895 0.315 1.785 ;
        RECT 3.610 1.625 3.780 1.785 ;
        RECT 3.610 1.455 5.205 1.625 ;
        RECT 5.035 1.245 5.205 1.455 ;
        RECT 5.035 1.075 5.745 1.245 ;
        RECT 0.085 0.645 0.910 0.895 ;
        RECT 1.130 0.725 2.320 0.905 ;
        RECT 1.130 0.475 1.380 0.725 ;
        RECT 0.105 0.255 1.380 0.475 ;
        RECT 1.600 0.085 1.770 0.555 ;
        RECT 1.940 0.255 2.320 0.725 ;
        RECT 2.630 0.085 2.800 0.905 ;
        RECT 2.970 0.725 5.755 0.905 ;
        RECT 2.970 0.255 3.350 0.725 ;
        RECT 3.570 0.085 3.740 0.555 ;
        RECT 3.910 0.255 4.325 0.725 ;
        RECT 5.405 0.645 5.755 0.725 ;
        RECT 4.545 0.085 4.715 0.555 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 2.665 2.125 2.835 2.295 ;
        RECT 3.685 2.125 3.855 2.295 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
      LAYER met1 ;
        RECT 2.605 2.280 2.895 2.325 ;
        RECT 3.625 2.280 3.915 2.325 ;
        RECT 2.605 2.140 3.915 2.280 ;
        RECT 2.605 2.095 2.895 2.140 ;
        RECT 3.625 2.095 3.915 2.140 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xnor2_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__xnor2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__xnor2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.040 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.220000 ;
    PORT
      LAYER li1 ;
        RECT 2.375 1.075 5.930 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.220000 ;
    PORT
      LAYER li1 ;
        RECT 1.835 1.445 6.270 1.615 ;
        RECT 1.835 1.275 2.005 1.445 ;
        RECT 0.490 1.075 2.005 1.275 ;
        RECT 6.100 1.275 6.270 1.445 ;
        RECT 6.100 1.075 8.170 1.275 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.040 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.060 0.105 11.030 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 11.230 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.040 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.858500 ;
    PORT
      LAYER li1 ;
        RECT 8.730 2.045 9.060 2.465 ;
        RECT 6.750 1.785 9.060 2.045 ;
        RECT 8.730 1.665 9.060 1.785 ;
        RECT 9.710 1.665 9.960 2.465 ;
        RECT 10.610 1.665 10.940 2.465 ;
        RECT 8.730 1.445 10.940 1.665 ;
        RECT 10.705 0.905 10.940 1.445 ;
        RECT 9.150 0.655 10.940 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 11.040 2.805 ;
        RECT 0.085 1.615 0.460 2.465 ;
        RECT 0.680 1.835 0.930 2.635 ;
        RECT 1.150 2.005 1.400 2.465 ;
        RECT 1.620 2.175 1.870 2.635 ;
        RECT 2.090 2.005 2.340 2.465 ;
        RECT 2.560 2.175 2.810 2.635 ;
        RECT 3.030 2.005 3.280 2.465 ;
        RECT 3.500 2.175 3.750 2.635 ;
        RECT 3.970 2.005 4.220 2.465 ;
        RECT 1.150 1.785 4.220 2.005 ;
        RECT 4.425 2.005 4.740 2.465 ;
        RECT 4.960 2.175 5.210 2.635 ;
        RECT 5.430 2.005 5.680 2.465 ;
        RECT 5.900 2.175 6.150 2.635 ;
        RECT 6.370 2.215 8.540 2.465 ;
        RECT 6.370 2.005 6.580 2.215 ;
        RECT 4.425 1.785 6.580 2.005 ;
        RECT 9.240 1.835 9.490 2.635 ;
        RECT 10.180 1.835 10.430 2.635 ;
        RECT 1.150 1.615 1.400 1.785 ;
        RECT 0.085 1.445 1.400 1.615 ;
        RECT 6.490 1.445 8.560 1.615 ;
        RECT 0.085 0.905 0.320 1.445 ;
        RECT 8.390 1.275 8.560 1.445 ;
        RECT 8.390 1.075 10.535 1.275 ;
        RECT 0.085 0.645 1.910 0.905 ;
        RECT 2.130 0.725 4.260 0.905 ;
        RECT 2.130 0.475 2.380 0.725 ;
        RECT 0.170 0.255 2.380 0.475 ;
        RECT 2.600 0.085 2.770 0.555 ;
        RECT 2.940 0.255 3.320 0.725 ;
        RECT 3.540 0.085 3.710 0.555 ;
        RECT 3.880 0.255 4.260 0.725 ;
        RECT 4.430 0.085 4.700 0.905 ;
        RECT 4.870 0.735 8.980 0.905 ;
        RECT 4.870 0.725 8.170 0.735 ;
        RECT 4.870 0.255 5.250 0.725 ;
        RECT 5.470 0.085 5.640 0.555 ;
        RECT 5.810 0.255 6.190 0.725 ;
        RECT 6.410 0.085 6.580 0.555 ;
        RECT 6.750 0.255 7.130 0.725 ;
        RECT 7.350 0.085 7.520 0.555 ;
        RECT 7.690 0.255 8.070 0.725 ;
        RECT 8.290 0.085 8.460 0.555 ;
        RECT 8.730 0.475 8.980 0.735 ;
        RECT 8.730 0.305 10.940 0.475 ;
        RECT 0.000 -0.085 11.040 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 1.165 1.445 1.335 1.615 ;
        RECT 6.725 1.445 6.895 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
      LAYER met1 ;
        RECT 1.055 1.600 1.395 1.645 ;
        RECT 6.655 1.600 7.005 1.645 ;
        RECT 1.055 1.460 7.005 1.600 ;
        RECT 1.055 1.415 1.395 1.460 ;
        RECT 6.655 1.415 7.005 1.460 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xnor2_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__xnor3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__xnor3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.200 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.276000 ;
    PORT
      LAYER li1 ;
        RECT 7.495 1.075 8.215 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.735900 ;
    PORT
      LAYER li1 ;
        RECT 6.625 1.445 7.255 1.615 ;
        RECT 6.625 0.995 6.845 1.445 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.425400 ;
    PORT
      LAYER li1 ;
        RECT 1.715 1.075 2.330 1.325 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.200 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.005 7.155 1.015 ;
        RECT 0.005 0.115 9.175 1.005 ;
        RECT 0.005 0.105 1.035 0.115 ;
        RECT 3.475 0.105 4.525 0.115 ;
        RECT 6.730 0.105 9.175 0.115 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.390 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.200 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.472000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.440 0.365 2.465 ;
        RECT 0.085 0.350 0.345 1.440 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.200 2.805 ;
        RECT 0.535 2.215 0.920 2.635 ;
        RECT 1.100 2.235 2.670 2.405 ;
        RECT 3.425 2.235 3.755 2.635 ;
        RECT 4.190 2.275 7.485 2.445 ;
        RECT 7.915 2.275 8.595 2.635 ;
        RECT 1.100 2.045 1.320 2.235 ;
        RECT 4.190 2.065 4.360 2.275 ;
        RECT 0.535 1.875 1.320 2.045 ;
        RECT 1.660 1.895 4.360 2.065 ;
        RECT 0.535 1.330 0.755 1.875 ;
        RECT 0.985 1.535 2.670 1.705 ;
        RECT 0.515 0.865 0.755 1.330 ;
        RECT 0.515 0.695 1.205 0.865 ;
        RECT 0.515 0.085 0.815 0.525 ;
        RECT 0.985 0.425 1.205 0.695 ;
        RECT 1.375 0.595 1.545 1.535 ;
        RECT 2.500 1.325 2.670 1.535 ;
        RECT 2.890 1.525 3.275 1.695 ;
        RECT 2.995 1.375 3.275 1.525 ;
        RECT 2.500 0.995 2.825 1.325 ;
        RECT 1.845 0.795 2.225 0.905 ;
        RECT 2.995 0.795 3.165 1.375 ;
        RECT 3.445 1.205 3.615 1.895 ;
        RECT 3.845 1.445 4.365 1.715 ;
        RECT 1.845 0.625 3.165 0.795 ;
        RECT 3.335 1.035 3.615 1.205 ;
        RECT 3.335 0.455 3.505 1.035 ;
        RECT 2.170 0.425 2.655 0.455 ;
        RECT 0.985 0.255 2.655 0.425 ;
        RECT 2.875 0.285 3.505 0.455 ;
        RECT 3.675 0.085 3.845 0.865 ;
        RECT 4.075 0.415 4.365 1.445 ;
        RECT 4.545 0.595 4.715 2.105 ;
        RECT 4.885 0.890 5.055 2.275 ;
        RECT 8.815 2.105 9.110 2.465 ;
        RECT 5.285 1.615 5.700 2.045 ;
        RECT 6.285 1.935 9.110 2.105 ;
        RECT 5.285 1.445 6.115 1.615 ;
        RECT 5.300 0.995 5.725 1.270 ;
        RECT 4.885 0.825 5.145 0.890 ;
        RECT 4.885 0.720 5.345 0.825 ;
        RECT 4.925 0.655 5.345 0.720 ;
        RECT 4.545 0.485 4.755 0.595 ;
        RECT 4.545 0.265 4.955 0.485 ;
        RECT 5.175 0.320 5.345 0.655 ;
        RECT 5.515 0.630 5.725 0.995 ;
        RECT 5.945 0.425 6.115 1.445 ;
        RECT 6.285 0.595 6.455 1.935 ;
        RECT 8.575 1.875 9.110 1.935 ;
        RECT 7.475 1.495 8.660 1.705 ;
        RECT 8.490 1.325 8.660 1.495 ;
        RECT 7.015 0.945 7.325 1.275 ;
        RECT 8.490 0.995 8.770 1.325 ;
        RECT 7.015 0.730 7.220 0.945 ;
        RECT 8.490 0.905 8.660 0.995 ;
        RECT 7.555 0.750 8.660 0.905 ;
        RECT 7.515 0.735 8.660 0.750 ;
        RECT 6.625 0.425 7.140 0.465 ;
        RECT 5.945 0.255 7.140 0.425 ;
        RECT 7.515 0.295 7.805 0.735 ;
        RECT 8.940 0.585 9.110 1.875 ;
        RECT 8.050 0.085 8.510 0.565 ;
        RECT 8.810 0.255 9.110 0.585 ;
        RECT 0.000 -0.085 9.200 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 3.105 1.445 3.275 1.615 ;
        RECT 4.075 0.765 4.245 0.935 ;
        RECT 5.555 1.445 5.725 1.615 ;
        RECT 4.585 0.425 4.755 0.595 ;
        RECT 5.555 0.765 5.725 0.935 ;
        RECT 7.035 0.765 7.205 0.935 ;
        RECT 7.545 0.425 7.715 0.595 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
      LAYER met1 ;
        RECT 3.045 1.600 3.335 1.645 ;
        RECT 5.495 1.600 5.785 1.645 ;
        RECT 3.045 1.460 5.785 1.600 ;
        RECT 3.045 1.415 3.335 1.460 ;
        RECT 5.495 1.415 5.785 1.460 ;
        RECT 4.015 0.920 4.305 0.965 ;
        RECT 5.495 0.920 5.785 0.965 ;
        RECT 6.975 0.920 7.265 0.965 ;
        RECT 4.015 0.780 7.265 0.920 ;
        RECT 4.015 0.735 4.305 0.780 ;
        RECT 5.495 0.735 5.785 0.780 ;
        RECT 6.975 0.735 7.265 0.780 ;
        RECT 4.525 0.580 4.815 0.625 ;
        RECT 7.485 0.580 7.775 0.625 ;
        RECT 4.525 0.440 7.775 0.580 ;
        RECT 4.525 0.395 4.815 0.440 ;
        RECT 7.485 0.395 7.775 0.440 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xnor3_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__xnor3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__xnor3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.660 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.276000 ;
    PORT
      LAYER li1 ;
        RECT 8.055 1.075 8.695 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.735900 ;
    PORT
      LAYER li1 ;
        RECT 7.135 1.445 7.765 1.615 ;
        RECT 7.135 0.995 7.355 1.445 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.425400 ;
    PORT
      LAYER li1 ;
        RECT 2.225 1.075 2.840 1.325 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.660 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.005 7.665 1.015 ;
        RECT 0.005 0.115 9.550 1.005 ;
        RECT 0.005 0.105 1.545 0.115 ;
        RECT 3.985 0.105 5.035 0.115 ;
        RECT 7.240 0.105 9.550 0.115 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.850 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.660 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.550500 ;
    PORT
      LAYER li1 ;
        RECT 0.545 0.350 0.865 2.465 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.660 2.805 ;
        RECT 0.085 1.490 0.375 2.635 ;
        RECT 1.045 2.215 1.430 2.635 ;
        RECT 1.610 2.235 3.180 2.405 ;
        RECT 3.935 2.235 4.265 2.635 ;
        RECT 4.700 2.275 7.995 2.445 ;
        RECT 8.455 2.275 8.790 2.635 ;
        RECT 1.610 2.045 1.830 2.235 ;
        RECT 4.700 2.065 4.870 2.275 ;
        RECT 1.045 1.875 1.830 2.045 ;
        RECT 2.170 1.895 4.870 2.065 ;
        RECT 1.045 0.865 1.265 1.875 ;
        RECT 1.495 1.535 3.180 1.705 ;
        RECT 0.085 0.085 0.375 0.735 ;
        RECT 1.045 0.695 1.715 0.865 ;
        RECT 1.035 0.085 1.325 0.525 ;
        RECT 1.495 0.425 1.715 0.695 ;
        RECT 1.885 0.595 2.055 1.535 ;
        RECT 3.010 1.325 3.180 1.535 ;
        RECT 3.400 1.525 3.785 1.695 ;
        RECT 3.505 1.375 3.785 1.525 ;
        RECT 3.010 0.995 3.335 1.325 ;
        RECT 2.355 0.795 2.735 0.905 ;
        RECT 3.505 0.795 3.675 1.375 ;
        RECT 3.955 1.205 4.125 1.895 ;
        RECT 4.355 1.445 4.875 1.715 ;
        RECT 2.355 0.625 3.675 0.795 ;
        RECT 3.845 1.035 4.125 1.205 ;
        RECT 3.845 0.455 4.015 1.035 ;
        RECT 2.680 0.425 3.165 0.455 ;
        RECT 1.495 0.255 3.165 0.425 ;
        RECT 3.385 0.285 4.015 0.455 ;
        RECT 4.185 0.085 4.355 0.865 ;
        RECT 4.585 0.415 4.875 1.445 ;
        RECT 5.055 0.595 5.225 2.105 ;
        RECT 5.395 0.890 5.565 2.275 ;
        RECT 9.190 2.105 9.485 2.465 ;
        RECT 5.795 1.615 6.210 2.045 ;
        RECT 6.795 1.935 9.485 2.105 ;
        RECT 5.795 1.445 6.625 1.615 ;
        RECT 5.810 0.995 6.235 1.270 ;
        RECT 5.395 0.825 5.655 0.890 ;
        RECT 5.395 0.720 5.855 0.825 ;
        RECT 5.435 0.655 5.855 0.720 ;
        RECT 5.055 0.485 5.265 0.595 ;
        RECT 5.055 0.265 5.465 0.485 ;
        RECT 5.685 0.320 5.855 0.655 ;
        RECT 6.025 0.630 6.235 0.995 ;
        RECT 6.455 0.425 6.625 1.445 ;
        RECT 6.795 0.595 6.965 1.935 ;
        RECT 8.950 1.875 9.485 1.935 ;
        RECT 7.985 1.495 9.035 1.705 ;
        RECT 8.865 1.325 9.035 1.495 ;
        RECT 7.525 0.945 7.835 1.275 ;
        RECT 8.865 0.995 9.145 1.325 ;
        RECT 7.525 0.730 7.730 0.945 ;
        RECT 8.865 0.905 9.035 0.995 ;
        RECT 8.065 0.750 9.035 0.905 ;
        RECT 8.025 0.735 9.035 0.750 ;
        RECT 7.135 0.425 7.650 0.465 ;
        RECT 6.455 0.255 7.650 0.425 ;
        RECT 8.025 0.295 8.315 0.735 ;
        RECT 9.315 0.585 9.485 1.875 ;
        RECT 8.535 0.085 8.705 0.565 ;
        RECT 9.185 0.255 9.485 0.585 ;
        RECT 0.000 -0.085 9.660 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 3.615 1.445 3.785 1.615 ;
        RECT 4.585 0.765 4.755 0.935 ;
        RECT 6.065 1.445 6.235 1.615 ;
        RECT 5.095 0.425 5.265 0.595 ;
        RECT 6.065 0.765 6.235 0.935 ;
        RECT 7.545 0.765 7.715 0.935 ;
        RECT 8.055 0.425 8.225 0.595 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
      LAYER met1 ;
        RECT 3.555 1.600 3.845 1.645 ;
        RECT 6.005 1.600 6.295 1.645 ;
        RECT 3.555 1.460 6.295 1.600 ;
        RECT 3.555 1.415 3.845 1.460 ;
        RECT 6.005 1.415 6.295 1.460 ;
        RECT 4.525 0.920 4.815 0.965 ;
        RECT 6.005 0.920 6.295 0.965 ;
        RECT 7.485 0.920 7.775 0.965 ;
        RECT 4.525 0.780 7.775 0.920 ;
        RECT 4.525 0.735 4.815 0.780 ;
        RECT 6.005 0.735 6.295 0.780 ;
        RECT 7.485 0.735 7.775 0.780 ;
        RECT 5.035 0.580 5.325 0.625 ;
        RECT 7.995 0.580 8.285 0.625 ;
        RECT 5.035 0.440 8.285 0.580 ;
        RECT 5.035 0.395 5.325 0.440 ;
        RECT 7.995 0.395 8.285 0.440 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xnor3_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__xnor3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__xnor3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.580 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.276000 ;
    PORT
      LAYER li1 ;
        RECT 9.075 1.075 9.535 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.735900 ;
    PORT
      LAYER li1 ;
        RECT 8.155 1.445 8.785 1.615 ;
        RECT 8.155 0.995 8.375 1.445 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.425400 ;
    PORT
      LAYER li1 ;
        RECT 3.245 1.075 3.860 1.325 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.580 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.115 1.005 8.685 1.015 ;
        RECT 0.115 0.115 10.390 1.005 ;
        RECT 0.115 0.105 2.565 0.115 ;
        RECT 5.005 0.105 6.065 0.115 ;
        RECT 8.260 0.105 10.390 0.115 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.770 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.580 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.996000 ;
    PORT
      LAYER li1 ;
        RECT 0.625 1.325 1.005 2.425 ;
        RECT 1.565 1.440 1.895 2.465 ;
        RECT 1.565 1.325 1.860 1.440 ;
        RECT 0.625 0.995 1.860 1.325 ;
        RECT 0.625 0.375 0.925 0.995 ;
        RECT 1.565 0.925 1.860 0.995 ;
        RECT 1.565 0.350 1.875 0.925 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.580 2.805 ;
        RECT 0.285 1.490 0.455 2.635 ;
        RECT 1.225 1.495 1.395 2.635 ;
        RECT 2.065 2.215 2.450 2.635 ;
        RECT 2.630 2.235 4.200 2.405 ;
        RECT 4.955 2.235 5.285 2.635 ;
        RECT 5.720 2.275 9.015 2.445 ;
        RECT 9.425 2.275 9.810 2.635 ;
        RECT 2.630 2.045 2.850 2.235 ;
        RECT 5.720 2.065 5.890 2.275 ;
        RECT 2.065 1.875 2.850 2.045 ;
        RECT 3.190 1.895 5.890 2.065 ;
        RECT 2.065 1.325 2.285 1.875 ;
        RECT 2.515 1.535 4.200 1.705 ;
        RECT 2.030 0.995 2.285 1.325 ;
        RECT 2.060 0.865 2.285 0.995 ;
        RECT 0.285 0.085 0.455 0.735 ;
        RECT 1.225 0.085 1.395 0.735 ;
        RECT 2.060 0.695 2.735 0.865 ;
        RECT 2.045 0.085 2.345 0.525 ;
        RECT 2.515 0.425 2.735 0.695 ;
        RECT 2.905 0.595 3.075 1.535 ;
        RECT 4.030 1.325 4.200 1.535 ;
        RECT 4.420 1.525 4.805 1.695 ;
        RECT 4.525 1.375 4.805 1.525 ;
        RECT 4.030 0.995 4.355 1.325 ;
        RECT 3.375 0.795 3.755 0.905 ;
        RECT 4.525 0.795 4.695 1.375 ;
        RECT 4.975 1.205 5.145 1.895 ;
        RECT 5.375 1.445 5.895 1.715 ;
        RECT 3.375 0.625 4.695 0.795 ;
        RECT 4.865 1.035 5.145 1.205 ;
        RECT 4.865 0.455 5.035 1.035 ;
        RECT 3.700 0.425 4.185 0.455 ;
        RECT 2.515 0.255 4.185 0.425 ;
        RECT 4.405 0.285 5.035 0.455 ;
        RECT 5.205 0.085 5.375 0.865 ;
        RECT 5.605 0.415 5.895 1.445 ;
        RECT 6.075 0.485 6.245 2.105 ;
        RECT 6.415 0.825 6.585 2.275 ;
        RECT 10.030 2.105 10.325 2.465 ;
        RECT 6.815 1.615 7.230 2.045 ;
        RECT 7.815 1.935 10.325 2.105 ;
        RECT 6.815 1.445 7.645 1.615 ;
        RECT 6.830 0.995 7.255 1.270 ;
        RECT 6.415 0.655 6.875 0.825 ;
        RECT 6.075 0.265 6.520 0.485 ;
        RECT 6.705 0.320 6.875 0.655 ;
        RECT 7.045 0.630 7.255 0.995 ;
        RECT 7.475 0.425 7.645 1.445 ;
        RECT 7.815 0.595 7.985 1.935 ;
        RECT 9.790 1.875 10.325 1.935 ;
        RECT 9.005 1.495 9.875 1.705 ;
        RECT 9.705 1.325 9.875 1.495 ;
        RECT 8.545 0.945 8.855 1.275 ;
        RECT 9.705 0.995 9.985 1.325 ;
        RECT 8.545 0.730 8.750 0.945 ;
        RECT 9.705 0.905 9.875 0.995 ;
        RECT 9.085 0.750 9.875 0.905 ;
        RECT 9.045 0.735 9.875 0.750 ;
        RECT 8.155 0.425 8.670 0.465 ;
        RECT 7.475 0.255 8.670 0.425 ;
        RECT 9.045 0.295 9.335 0.735 ;
        RECT 10.155 0.585 10.325 1.875 ;
        RECT 9.555 0.085 9.725 0.565 ;
        RECT 10.025 0.255 10.325 0.585 ;
        RECT 0.000 -0.085 10.580 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 4.635 1.445 4.805 1.615 ;
        RECT 5.605 0.765 5.775 0.935 ;
        RECT 7.085 1.445 7.255 1.615 ;
        RECT 6.075 0.425 6.245 0.595 ;
        RECT 7.085 0.765 7.255 0.935 ;
        RECT 8.565 0.765 8.735 0.935 ;
        RECT 9.075 0.425 9.245 0.595 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
      LAYER met1 ;
        RECT 4.575 1.600 4.865 1.645 ;
        RECT 7.025 1.600 7.315 1.645 ;
        RECT 4.575 1.460 7.315 1.600 ;
        RECT 4.575 1.415 4.865 1.460 ;
        RECT 7.025 1.415 7.315 1.460 ;
        RECT 5.545 0.920 5.835 0.965 ;
        RECT 7.025 0.920 7.315 0.965 ;
        RECT 8.505 0.920 8.795 0.965 ;
        RECT 5.545 0.780 8.795 0.920 ;
        RECT 5.545 0.735 5.835 0.780 ;
        RECT 7.025 0.735 7.315 0.780 ;
        RECT 8.505 0.735 8.795 0.780 ;
        RECT 6.015 0.580 6.315 0.625 ;
        RECT 9.015 0.580 9.305 0.625 ;
        RECT 6.015 0.440 9.305 0.580 ;
        RECT 6.015 0.395 6.315 0.440 ;
        RECT 9.015 0.395 9.305 0.440 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xnor3_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__xor2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__xor2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.955 1.075 1.500 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.555000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.445 1.890 1.615 ;
        RECT 0.425 0.995 0.775 1.445 ;
        RECT 1.720 1.245 1.890 1.445 ;
        RECT 1.720 1.075 2.155 1.245 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.045 0.105 3.625 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.996000 ;
    PORT
      LAYER li1 ;
        RECT 3.225 1.535 3.545 2.465 ;
        RECT 2.915 1.365 3.545 1.535 ;
        RECT 2.915 0.485 3.085 1.365 ;
        RECT 1.880 0.315 3.085 0.485 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.085 1.785 0.465 2.465 ;
        RECT 1.165 1.785 1.335 2.635 ;
        RECT 1.505 1.955 1.885 2.465 ;
        RECT 2.115 2.125 2.285 2.635 ;
        RECT 2.455 1.955 2.855 2.465 ;
        RECT 1.505 1.785 2.855 1.955 ;
        RECT 0.085 0.825 0.255 1.785 ;
        RECT 2.515 0.825 2.745 1.325 ;
        RECT 0.085 0.655 2.745 0.825 ;
        RECT 0.135 0.085 0.465 0.475 ;
        RECT 0.685 0.335 0.855 0.655 ;
        RECT 1.035 0.085 1.415 0.475 ;
        RECT 3.255 0.085 3.545 0.920 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xor2_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__xor2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__xor2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER li1 ;
        RECT 0.755 1.445 2.080 1.615 ;
        RECT 0.755 1.275 0.925 1.445 ;
        RECT 0.545 1.075 0.925 1.275 ;
        RECT 1.860 1.275 2.080 1.445 ;
        RECT 1.860 1.075 3.530 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER met1 ;
        RECT 1.105 1.260 1.395 1.305 ;
        RECT 3.765 1.260 4.055 1.305 ;
        RECT 1.105 1.120 4.055 1.260 ;
        RECT 1.105 1.075 1.395 1.120 ;
        RECT 3.765 1.075 4.055 1.120 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 6.325 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.806750 ;
    PORT
      LAYER li1 ;
        RECT 5.475 1.625 5.725 2.125 ;
        RECT 5.475 1.415 6.350 1.625 ;
        RECT 5.985 0.905 6.350 1.415 ;
        RECT 3.975 0.725 6.350 0.905 ;
        RECT 3.975 0.645 4.305 0.725 ;
        RECT 5.385 0.645 5.765 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.120 2.135 0.400 2.465 ;
        RECT 0.620 2.135 0.870 2.635 ;
        RECT 1.090 2.295 2.280 2.465 ;
        RECT 1.090 2.135 1.340 2.295 ;
        RECT 2.030 2.135 2.280 2.295 ;
        RECT 0.145 2.125 0.315 2.135 ;
        RECT 1.165 2.125 1.335 2.135 ;
        RECT 2.485 2.125 2.800 2.465 ;
        RECT 3.020 2.135 3.270 2.635 ;
        RECT 1.560 1.955 1.810 2.125 ;
        RECT 2.590 1.955 2.800 2.125 ;
        RECT 3.490 1.955 3.740 2.465 ;
        RECT 3.960 2.135 4.265 2.635 ;
        RECT 4.485 2.295 6.195 2.465 ;
        RECT 4.485 1.955 5.255 2.295 ;
        RECT 0.120 1.785 2.420 1.955 ;
        RECT 2.590 1.785 5.255 1.955 ;
        RECT 5.945 1.795 6.195 2.295 ;
        RECT 0.120 0.905 0.290 1.785 ;
        RECT 2.250 1.615 2.420 1.785 ;
        RECT 2.250 1.445 5.185 1.615 ;
        RECT 1.145 1.075 1.690 1.275 ;
        RECT 3.720 1.075 4.490 1.275 ;
        RECT 5.015 1.245 5.185 1.445 ;
        RECT 5.015 1.075 5.725 1.245 ;
        RECT 0.120 0.725 1.850 0.905 ;
        RECT 0.190 0.085 0.360 0.555 ;
        RECT 0.530 0.255 0.910 0.725 ;
        RECT 1.130 0.085 1.300 0.555 ;
        RECT 1.470 0.255 1.850 0.725 ;
        RECT 2.510 0.725 3.700 0.905 ;
        RECT 2.070 0.085 2.240 0.555 ;
        RECT 2.510 0.255 2.840 0.725 ;
        RECT 3.060 0.085 3.230 0.555 ;
        RECT 3.400 0.475 3.700 0.725 ;
        RECT 3.400 0.255 4.780 0.475 ;
        RECT 5.045 0.085 5.215 0.555 ;
        RECT 5.985 0.085 6.155 0.555 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 1.165 1.105 1.335 1.275 ;
        RECT 3.825 1.105 3.995 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
      LAYER met1 ;
        RECT 0.085 2.280 0.375 2.325 ;
        RECT 1.105 2.280 1.395 2.325 ;
        RECT 0.085 2.140 1.395 2.280 ;
        RECT 0.085 2.095 0.375 2.140 ;
        RECT 1.105 2.095 1.395 2.140 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xor2_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__xor2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__xor2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.040 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.220000 ;
    PORT
      LAYER li1 ;
        RECT 2.880 1.445 6.815 1.615 ;
        RECT 2.880 1.275 3.100 1.445 ;
        RECT 0.425 1.075 3.100 1.275 ;
        RECT 6.595 1.275 6.815 1.445 ;
        RECT 6.595 1.075 8.120 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.220000 ;
    PORT
      LAYER li1 ;
        RECT 3.270 1.105 6.340 1.275 ;
        RECT 3.270 1.075 5.500 1.105 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.040 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 11.000 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 11.230 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.040 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.759450 ;
    PORT
      LAYER met1 ;
        RECT 5.645 0.780 8.995 0.925 ;
        RECT 5.645 0.695 5.935 0.780 ;
        RECT 8.705 0.695 8.995 0.780 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 11.040 2.805 ;
        RECT 0.085 2.005 0.400 2.465 ;
        RECT 0.620 2.175 0.870 2.635 ;
        RECT 1.090 2.005 1.340 2.465 ;
        RECT 1.560 2.175 1.810 2.635 ;
        RECT 2.030 2.295 4.160 2.465 ;
        RECT 2.030 2.005 2.280 2.295 ;
        RECT 2.970 2.125 3.220 2.295 ;
        RECT 0.085 1.785 2.280 2.005 ;
        RECT 2.500 1.955 2.750 2.125 ;
        RECT 3.440 1.955 3.690 2.125 ;
        RECT 2.500 1.785 3.690 1.955 ;
        RECT 3.910 1.795 4.160 2.295 ;
        RECT 4.430 2.005 4.680 2.465 ;
        RECT 4.900 2.175 5.150 2.635 ;
        RECT 5.370 2.005 5.620 2.465 ;
        RECT 5.840 2.175 6.090 2.635 ;
        RECT 6.310 2.005 6.560 2.465 ;
        RECT 6.780 2.175 7.030 2.635 ;
        RECT 7.250 2.005 7.500 2.465 ;
        RECT 7.720 2.175 7.970 2.635 ;
        RECT 8.190 2.295 10.380 2.465 ;
        RECT 8.190 2.005 8.440 2.295 ;
        RECT 4.430 1.785 8.440 2.005 ;
        RECT 2.500 1.615 2.670 1.785 ;
        RECT 0.085 1.445 2.670 1.615 ;
        RECT 7.250 1.455 7.500 1.785 ;
        RECT 8.680 1.665 8.970 2.125 ;
        RECT 9.190 1.835 9.440 2.295 ;
        RECT 9.660 1.665 9.910 2.125 ;
        RECT 10.130 1.795 10.380 2.295 ;
        RECT 8.680 1.625 9.910 1.665 ;
        RECT 10.550 1.625 10.955 2.465 ;
        RECT 8.010 1.445 8.510 1.615 ;
        RECT 8.680 1.445 10.955 1.625 ;
        RECT 0.085 0.905 0.255 1.445 ;
        RECT 8.340 1.275 8.510 1.445 ;
        RECT 8.340 1.075 10.130 1.275 ;
        RECT 5.650 0.905 6.130 0.935 ;
        RECT 10.635 0.905 10.955 1.445 ;
        RECT 0.085 0.735 3.730 0.905 ;
        RECT 0.530 0.725 3.730 0.735 ;
        RECT 0.085 0.085 0.360 0.565 ;
        RECT 0.530 0.255 0.910 0.725 ;
        RECT 1.130 0.085 1.300 0.555 ;
        RECT 1.470 0.255 1.850 0.725 ;
        RECT 2.070 0.085 2.240 0.555 ;
        RECT 2.410 0.255 2.790 0.725 ;
        RECT 3.010 0.085 3.180 0.555 ;
        RECT 3.350 0.255 3.730 0.725 ;
        RECT 3.950 0.085 4.220 0.895 ;
        RECT 4.565 0.645 6.130 0.905 ;
        RECT 6.350 0.725 8.480 0.905 ;
        RECT 8.650 0.735 10.955 0.905 ;
        RECT 8.650 0.725 9.480 0.735 ;
        RECT 6.350 0.475 6.600 0.725 ;
        RECT 4.390 0.255 6.600 0.475 ;
        RECT 6.820 0.085 6.990 0.555 ;
        RECT 7.160 0.255 7.540 0.725 ;
        RECT 7.760 0.085 7.930 0.555 ;
        RECT 8.100 0.255 8.480 0.725 ;
        RECT 8.760 0.085 8.930 0.555 ;
        RECT 9.100 0.255 9.480 0.725 ;
        RECT 9.700 0.085 9.870 0.555 ;
        RECT 10.040 0.255 10.420 0.735 ;
        RECT 10.640 0.085 10.810 0.555 ;
        RECT 0.000 -0.085 11.040 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 2.185 1.445 2.355 1.615 ;
        RECT 8.305 1.445 8.475 1.615 ;
        RECT 5.705 0.725 5.875 0.895 ;
        RECT 8.765 0.725 8.935 0.895 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
      LAYER met1 ;
        RECT 2.125 1.600 2.415 1.645 ;
        RECT 8.245 1.600 8.535 1.645 ;
        RECT 2.125 1.460 8.535 1.600 ;
        RECT 2.125 1.415 2.415 1.460 ;
        RECT 8.245 1.415 8.535 1.460 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xor2_4

#--------EOF---------

MACRO sky130_fd_sc_hdll__xor3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__xor3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.660 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.276000 ;
    PORT
      LAYER li1 ;
        RECT 8.005 1.075 8.695 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.735900 ;
    PORT
      LAYER li1 ;
        RECT 7.085 1.445 7.715 1.725 ;
        RECT 7.085 0.995 7.305 1.445 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.425400 ;
    PORT
      LAYER li1 ;
        RECT 1.960 0.995 2.645 1.325 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.660 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.170 1.005 7.615 1.015 ;
        RECT 0.170 0.115 9.630 1.005 ;
        RECT 0.170 0.105 1.285 0.115 ;
        RECT 3.920 0.105 4.980 0.115 ;
        RECT 7.190 0.105 9.630 0.115 ;
        RECT 0.170 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.850 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.660 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.472000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.440 0.610 2.465 ;
        RECT 0.085 0.925 0.400 1.440 ;
        RECT 0.085 0.350 0.590 0.925 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.660 2.805 ;
        RECT 0.830 2.215 1.165 2.635 ;
        RECT 1.350 2.235 3.045 2.405 ;
        RECT 3.310 2.235 3.715 2.405 ;
        RECT 3.885 2.235 4.215 2.635 ;
        RECT 4.650 2.275 7.945 2.445 ;
        RECT 8.355 2.275 9.050 2.635 ;
        RECT 1.350 2.045 1.570 2.235 ;
        RECT 3.545 2.065 3.715 2.235 ;
        RECT 4.650 2.065 4.820 2.275 ;
        RECT 0.800 1.875 1.570 2.045 ;
        RECT 1.970 1.895 3.375 2.065 ;
        RECT 3.545 1.895 4.820 2.065 ;
        RECT 0.800 0.865 1.000 1.875 ;
        RECT 1.235 1.535 2.985 1.705 ;
        RECT 0.800 0.695 1.450 0.865 ;
        RECT 0.810 0.085 1.060 0.525 ;
        RECT 1.230 0.425 1.450 0.695 ;
        RECT 1.620 0.595 1.790 1.535 ;
        RECT 2.815 1.325 2.985 1.535 ;
        RECT 3.205 1.695 3.375 1.895 ;
        RECT 3.205 1.525 3.735 1.695 ;
        RECT 3.450 1.375 3.735 1.525 ;
        RECT 2.815 0.995 3.140 1.325 ;
        RECT 2.070 0.655 3.280 0.825 ;
        RECT 2.490 0.425 2.890 0.455 ;
        RECT 1.230 0.255 2.890 0.425 ;
        RECT 3.060 0.425 3.280 0.655 ;
        RECT 3.450 0.595 3.620 1.375 ;
        RECT 3.905 1.205 4.075 1.895 ;
        RECT 4.305 1.445 4.820 1.715 ;
        RECT 3.790 1.035 4.075 1.205 ;
        RECT 3.790 0.425 3.960 1.035 ;
        RECT 3.060 0.255 3.960 0.425 ;
        RECT 4.130 0.085 4.300 0.865 ;
        RECT 4.530 0.415 4.820 1.445 ;
        RECT 4.995 0.595 5.165 2.105 ;
        RECT 5.335 0.890 5.505 2.275 ;
        RECT 9.270 2.105 9.565 2.465 ;
        RECT 5.745 1.615 6.160 2.045 ;
        RECT 6.745 1.935 9.565 2.105 ;
        RECT 5.745 1.445 6.575 1.615 ;
        RECT 5.760 0.995 6.185 1.270 ;
        RECT 5.335 0.825 5.605 0.890 ;
        RECT 5.335 0.720 5.800 0.825 ;
        RECT 5.385 0.655 5.800 0.720 ;
        RECT 4.995 0.485 5.215 0.595 ;
        RECT 4.995 0.265 5.410 0.485 ;
        RECT 5.630 0.320 5.800 0.655 ;
        RECT 5.970 0.630 6.185 0.995 ;
        RECT 6.405 0.425 6.575 1.445 ;
        RECT 6.745 0.595 6.915 1.935 ;
        RECT 9.030 1.875 9.565 1.935 ;
        RECT 7.935 1.495 9.115 1.705 ;
        RECT 8.945 1.325 9.115 1.495 ;
        RECT 7.475 0.945 7.785 1.275 ;
        RECT 8.945 0.995 9.225 1.325 ;
        RECT 7.475 0.730 7.680 0.945 ;
        RECT 8.945 0.905 9.115 0.995 ;
        RECT 8.015 0.750 9.115 0.905 ;
        RECT 7.975 0.735 9.115 0.750 ;
        RECT 7.085 0.425 7.600 0.465 ;
        RECT 6.405 0.255 7.600 0.425 ;
        RECT 7.975 0.295 8.265 0.735 ;
        RECT 9.395 0.585 9.565 1.875 ;
        RECT 8.485 0.085 8.935 0.565 ;
        RECT 9.265 0.255 9.565 0.585 ;
        RECT 0.000 -0.085 9.660 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 3.565 1.445 3.735 1.615 ;
        RECT 4.535 0.765 4.705 0.935 ;
        RECT 6.015 1.445 6.185 1.615 ;
        RECT 5.045 0.425 5.215 0.595 ;
        RECT 6.015 0.765 6.185 0.935 ;
        RECT 7.495 0.765 7.665 0.935 ;
        RECT 8.005 0.425 8.175 0.595 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
      LAYER met1 ;
        RECT 3.505 1.600 3.795 1.645 ;
        RECT 5.955 1.600 6.245 1.645 ;
        RECT 3.505 1.460 6.245 1.600 ;
        RECT 3.505 1.415 3.795 1.460 ;
        RECT 5.955 1.415 6.245 1.460 ;
        RECT 4.475 0.920 4.765 0.965 ;
        RECT 5.955 0.920 6.245 0.965 ;
        RECT 7.435 0.920 7.725 0.965 ;
        RECT 4.475 0.780 7.725 0.920 ;
        RECT 4.475 0.735 4.765 0.780 ;
        RECT 5.955 0.735 6.245 0.780 ;
        RECT 7.435 0.735 7.725 0.780 ;
        RECT 4.985 0.580 5.275 0.625 ;
        RECT 7.945 0.580 8.235 0.625 ;
        RECT 4.985 0.440 8.235 0.580 ;
        RECT 4.985 0.395 5.275 0.440 ;
        RECT 7.945 0.395 8.235 0.440 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xor3_1

#--------EOF---------

MACRO sky130_fd_sc_hdll__xor3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__xor3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.660 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.276000 ;
    PORT
      LAYER li1 ;
        RECT 8.300 1.075 8.760 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.735900 ;
    PORT
      LAYER li1 ;
        RECT 7.380 1.445 8.010 1.665 ;
        RECT 7.380 0.995 7.600 1.445 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.425400 ;
    PORT
      LAYER li1 ;
        RECT 2.255 0.995 2.940 1.325 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.660 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.005 7.910 1.015 ;
        RECT 0.005 0.115 9.590 1.005 ;
        RECT 0.005 0.105 1.580 0.115 ;
        RECT 4.215 0.105 5.275 0.115 ;
        RECT 7.485 0.105 9.590 0.115 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.850 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.660 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.517500 ;
    PORT
      LAYER li1 ;
        RECT 0.655 2.045 0.905 2.465 ;
        RECT 0.330 1.440 0.905 2.045 ;
        RECT 0.330 0.925 0.695 1.440 ;
        RECT 0.330 0.660 0.930 0.925 ;
        RECT 0.680 0.350 0.930 0.660 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.660 2.805 ;
        RECT 0.105 2.215 0.435 2.635 ;
        RECT 1.125 2.215 1.460 2.635 ;
        RECT 1.645 2.235 3.340 2.405 ;
        RECT 3.605 2.235 4.010 2.405 ;
        RECT 4.180 2.235 4.510 2.635 ;
        RECT 4.945 2.275 8.240 2.445 ;
        RECT 8.650 2.275 9.035 2.635 ;
        RECT 1.645 2.045 1.865 2.235 ;
        RECT 3.840 2.065 4.010 2.235 ;
        RECT 4.945 2.065 5.115 2.275 ;
        RECT 1.125 1.875 1.865 2.045 ;
        RECT 2.265 1.895 3.670 2.065 ;
        RECT 3.840 1.895 5.115 2.065 ;
        RECT 1.125 1.325 1.295 1.875 ;
        RECT 1.530 1.535 3.280 1.705 ;
        RECT 1.095 0.995 1.295 1.325 ;
        RECT 1.125 0.865 1.295 0.995 ;
        RECT 1.125 0.695 1.745 0.865 ;
        RECT 0.105 0.085 0.435 0.465 ;
        RECT 1.105 0.085 1.355 0.525 ;
        RECT 1.525 0.425 1.745 0.695 ;
        RECT 1.915 0.595 2.085 1.535 ;
        RECT 3.110 1.325 3.280 1.535 ;
        RECT 3.500 1.695 3.670 1.895 ;
        RECT 3.500 1.525 4.030 1.695 ;
        RECT 3.745 1.375 4.030 1.525 ;
        RECT 3.110 0.995 3.435 1.325 ;
        RECT 2.365 0.655 3.575 0.825 ;
        RECT 2.785 0.425 3.190 0.455 ;
        RECT 1.525 0.255 3.190 0.425 ;
        RECT 3.360 0.425 3.575 0.655 ;
        RECT 3.745 0.595 3.915 1.375 ;
        RECT 4.200 1.205 4.370 1.895 ;
        RECT 4.600 1.445 5.115 1.715 ;
        RECT 4.085 1.035 4.370 1.205 ;
        RECT 4.085 0.425 4.255 1.035 ;
        RECT 3.360 0.255 4.255 0.425 ;
        RECT 4.425 0.085 4.595 0.865 ;
        RECT 4.825 0.415 5.115 1.445 ;
        RECT 5.290 0.595 5.460 2.105 ;
        RECT 5.630 0.890 5.800 2.275 ;
        RECT 9.255 2.105 9.550 2.465 ;
        RECT 6.040 1.615 6.455 2.045 ;
        RECT 7.040 1.935 9.550 2.105 ;
        RECT 6.040 1.445 6.870 1.615 ;
        RECT 6.055 0.995 6.480 1.270 ;
        RECT 5.630 0.825 5.900 0.890 ;
        RECT 5.630 0.720 6.095 0.825 ;
        RECT 5.680 0.655 6.095 0.720 ;
        RECT 5.290 0.485 5.510 0.595 ;
        RECT 5.290 0.265 5.705 0.485 ;
        RECT 5.925 0.320 6.095 0.655 ;
        RECT 6.265 0.630 6.480 0.995 ;
        RECT 6.700 0.425 6.870 1.445 ;
        RECT 7.040 0.595 7.210 1.935 ;
        RECT 9.015 1.875 9.550 1.935 ;
        RECT 8.230 1.495 9.100 1.705 ;
        RECT 8.930 1.325 9.100 1.495 ;
        RECT 7.770 0.945 8.090 1.275 ;
        RECT 8.930 0.995 9.210 1.325 ;
        RECT 7.770 0.730 7.975 0.945 ;
        RECT 8.930 0.905 9.100 0.995 ;
        RECT 8.310 0.750 9.100 0.905 ;
        RECT 8.270 0.735 9.100 0.750 ;
        RECT 7.380 0.425 7.895 0.465 ;
        RECT 6.700 0.255 7.895 0.425 ;
        RECT 8.270 0.295 8.560 0.735 ;
        RECT 9.380 0.585 9.550 1.875 ;
        RECT 8.780 0.085 8.950 0.565 ;
        RECT 9.250 0.255 9.550 0.585 ;
        RECT 0.000 -0.085 9.660 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 3.860 1.445 4.030 1.615 ;
        RECT 4.830 0.765 5.000 0.935 ;
        RECT 6.310 1.445 6.480 1.615 ;
        RECT 5.340 0.425 5.510 0.595 ;
        RECT 6.310 0.765 6.480 0.935 ;
        RECT 7.790 0.765 7.960 0.935 ;
        RECT 8.300 0.425 8.470 0.595 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
      LAYER met1 ;
        RECT 3.800 1.600 4.090 1.645 ;
        RECT 6.250 1.600 6.540 1.645 ;
        RECT 3.800 1.460 6.540 1.600 ;
        RECT 3.800 1.415 4.090 1.460 ;
        RECT 6.250 1.415 6.540 1.460 ;
        RECT 4.770 0.920 5.060 0.965 ;
        RECT 6.250 0.920 6.540 0.965 ;
        RECT 7.730 0.920 8.020 0.965 ;
        RECT 4.770 0.780 8.020 0.920 ;
        RECT 4.770 0.735 5.060 0.780 ;
        RECT 6.250 0.735 6.540 0.780 ;
        RECT 7.730 0.735 8.020 0.780 ;
        RECT 5.280 0.580 5.570 0.625 ;
        RECT 8.240 0.580 8.530 0.625 ;
        RECT 5.280 0.440 8.530 0.580 ;
        RECT 5.280 0.395 5.570 0.440 ;
        RECT 8.240 0.395 8.530 0.440 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xor3_2

#--------EOF---------

MACRO sky130_fd_sc_hdll__xor3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__xor3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.580 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.276000 ;
    PORT
      LAYER li1 ;
        RECT 9.175 1.075 9.635 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.735900 ;
    PORT
      LAYER li1 ;
        RECT 8.255 1.445 8.640 1.615 ;
        RECT 8.255 0.995 8.475 1.445 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.425400 ;
    PORT
      LAYER li1 ;
        RECT 3.130 0.995 3.815 1.325 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.580 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.005 8.785 1.015 ;
        RECT 0.005 0.115 10.505 1.005 ;
        RECT 0.005 0.105 2.595 0.115 ;
        RECT 5.130 0.105 6.150 0.115 ;
        RECT 8.360 0.105 10.505 0.115 ;
        RECT 0.235 -0.085 0.405 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.770 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.580 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.996000 ;
    PORT
      LAYER li1 ;
        RECT 0.745 2.045 0.915 2.465 ;
        RECT 1.685 2.045 1.855 2.465 ;
        RECT 0.745 1.455 1.855 2.045 ;
        RECT 0.745 1.440 1.570 1.455 ;
        RECT 1.205 0.925 1.570 1.440 ;
        RECT 0.645 0.660 1.755 0.925 ;
        RECT 0.645 0.350 0.815 0.660 ;
        RECT 1.585 0.350 1.755 0.660 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.580 2.805 ;
        RECT 0.275 2.135 0.445 2.635 ;
        RECT 1.135 2.215 1.465 2.635 ;
        RECT 2.075 2.215 2.405 2.635 ;
        RECT 2.575 2.235 4.215 2.405 ;
        RECT 4.480 2.235 4.885 2.405 ;
        RECT 5.055 2.235 5.385 2.635 ;
        RECT 5.820 2.275 9.115 2.445 ;
        RECT 9.615 2.275 9.945 2.635 ;
        RECT 2.575 2.045 2.795 2.235 ;
        RECT 4.715 2.065 4.885 2.235 ;
        RECT 5.820 2.065 5.990 2.275 ;
        RECT 2.075 1.875 2.795 2.045 ;
        RECT 3.140 1.895 4.545 2.065 ;
        RECT 4.715 1.895 5.990 2.065 ;
        RECT 2.075 1.325 2.245 1.875 ;
        RECT 2.570 1.535 4.155 1.705 ;
        RECT 2.020 0.965 2.245 1.325 ;
        RECT 2.075 0.865 2.245 0.965 ;
        RECT 2.075 0.695 2.565 0.865 ;
        RECT 0.175 0.085 0.345 0.545 ;
        RECT 0.985 0.085 1.365 0.465 ;
        RECT 2.055 0.085 2.225 0.525 ;
        RECT 2.395 0.425 2.565 0.695 ;
        RECT 2.790 0.595 2.960 1.535 ;
        RECT 3.985 1.325 4.155 1.535 ;
        RECT 4.375 1.695 4.545 1.895 ;
        RECT 4.375 1.525 4.905 1.695 ;
        RECT 4.620 1.375 4.905 1.525 ;
        RECT 3.985 0.995 4.405 1.325 ;
        RECT 3.240 0.655 4.450 0.825 ;
        RECT 3.660 0.425 4.060 0.455 ;
        RECT 2.395 0.255 4.060 0.425 ;
        RECT 4.230 0.425 4.450 0.655 ;
        RECT 4.620 0.595 4.790 1.375 ;
        RECT 5.075 1.205 5.245 1.895 ;
        RECT 5.475 1.445 5.990 1.715 ;
        RECT 4.960 1.050 5.245 1.205 ;
        RECT 4.960 1.045 5.240 1.050 ;
        RECT 4.960 1.040 5.230 1.045 ;
        RECT 4.960 1.035 5.215 1.040 ;
        RECT 4.960 0.425 5.130 1.035 ;
        RECT 4.230 0.255 5.130 0.425 ;
        RECT 5.300 0.085 5.470 0.885 ;
        RECT 5.700 0.415 5.990 1.445 ;
        RECT 6.165 0.595 6.335 2.105 ;
        RECT 6.525 0.890 6.695 2.275 ;
        RECT 10.165 2.105 10.425 2.465 ;
        RECT 6.915 1.615 7.330 2.045 ;
        RECT 7.915 1.935 10.425 2.105 ;
        RECT 6.915 1.445 7.745 1.615 ;
        RECT 6.930 0.995 7.355 1.270 ;
        RECT 6.525 0.825 6.775 0.890 ;
        RECT 6.525 0.720 6.970 0.825 ;
        RECT 6.555 0.655 6.970 0.720 ;
        RECT 6.165 0.485 6.385 0.595 ;
        RECT 6.165 0.265 6.580 0.485 ;
        RECT 6.800 0.320 6.970 0.655 ;
        RECT 7.140 0.630 7.355 0.995 ;
        RECT 7.575 0.425 7.745 1.445 ;
        RECT 7.915 0.595 8.085 1.935 ;
        RECT 9.890 1.875 10.425 1.935 ;
        RECT 9.105 1.495 9.975 1.705 ;
        RECT 9.805 1.325 9.975 1.495 ;
        RECT 8.645 0.945 8.955 1.275 ;
        RECT 9.805 0.995 10.035 1.325 ;
        RECT 8.645 0.730 8.850 0.945 ;
        RECT 9.805 0.905 9.975 0.995 ;
        RECT 9.185 0.750 9.975 0.905 ;
        RECT 9.145 0.735 9.975 0.750 ;
        RECT 8.255 0.425 8.770 0.465 ;
        RECT 7.575 0.255 8.770 0.425 ;
        RECT 9.145 0.295 9.435 0.735 ;
        RECT 10.255 0.585 10.425 1.875 ;
        RECT 9.695 0.085 9.865 0.565 ;
        RECT 10.165 0.255 10.425 0.585 ;
        RECT 0.000 -0.085 10.580 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 4.735 1.445 4.905 1.615 ;
        RECT 5.705 0.765 5.875 0.935 ;
        RECT 7.185 1.445 7.355 1.615 ;
        RECT 6.215 0.425 6.385 0.595 ;
        RECT 7.185 0.765 7.355 0.935 ;
        RECT 8.665 0.765 8.835 0.935 ;
        RECT 9.175 0.425 9.345 0.595 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
      LAYER met1 ;
        RECT 4.675 1.600 4.965 1.645 ;
        RECT 7.125 1.600 7.415 1.645 ;
        RECT 4.675 1.460 7.415 1.600 ;
        RECT 4.675 1.415 4.965 1.460 ;
        RECT 7.125 1.415 7.415 1.460 ;
        RECT 5.645 0.920 5.985 0.965 ;
        RECT 7.125 0.920 7.415 0.965 ;
        RECT 8.605 0.920 8.895 0.965 ;
        RECT 5.645 0.780 8.895 0.920 ;
        RECT 5.645 0.735 5.985 0.780 ;
        RECT 7.125 0.735 7.415 0.780 ;
        RECT 8.605 0.735 8.895 0.780 ;
        RECT 6.155 0.580 6.445 0.625 ;
        RECT 9.115 0.580 9.405 0.625 ;
        RECT 6.155 0.440 9.405 0.580 ;
        RECT 6.155 0.395 6.445 0.440 ;
        RECT 9.115 0.395 9.405 0.440 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xor3_4

#--------EOF---------


END LIBRARY
