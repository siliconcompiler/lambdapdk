// //#############################################################################
// //# Function: Synchronizer with async reset                                   #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// module la_drsync
//   #(parameter PROP = "DEFAULT")
//    (
//     input  clk,    // clock
//     input  in,     // input data
//     input  nreset, // async active low reset
//     output out     // synchronized data
//     );
// 
//    localparam STAGES=2;
// 
//    reg [STAGES-1:0] shiftreg;
// 
//    always @ (posedge clk or negedge nreset)
//      if(!nreset)
//        shiftreg[STAGES-1:0] <= 'b0;
//      else
//        shiftreg[STAGES-1:0] <= {shiftreg[STAGES-2:0],in};
// 
//    assign out = shiftreg[STAGES-1];
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_drsync(clk, in, nreset, out);
  wire _0_;
  wire _1_;
  wire _2_;
  wire _3_;
  input clk;
  wire clk;
  input in;
  wire in;
  input nreset;
  wire nreset;
  output out;
  wire out;
  wire \shiftreg[0] ;
  INVx2_ASAP7_75t_R _4_ (
    .A(nreset),
    .Y(_2_)
  );
  INVx2_ASAP7_75t_R _5_ (
    .A(_0_),
    .Y(out)
  );
  INVx2_ASAP7_75t_R _6_ (
    .A(_1_),
    .Y(\shiftreg[0] )
  );
  ASYNC_DFFHx1_ASAP7_75t_R _7_ (
    .CLK(clk),
    .D(in),
    .QN(_1_),
    .RESET(_2_),
    .SET(_3_)
  );
  ASYNC_DFFHx1_ASAP7_75t_R _8_ (
    .CLK(clk),
    .D(\shiftreg[0] ),
    .QN(_0_),
    .RESET(_2_),
    .SET(_3_)
  );
  TIELOx1_ASAP7_75t_R _9_ (
    .L(_3_)
  );
endmodule
