VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram45_128x32
  FOREIGN fakeram45_128x32 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 78.470 BY 42.000 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.100 0.070 2.170 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.310 0.070 2.380 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.520 0.070 2.590 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.730 0.070 2.800 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.940 0.070 3.010 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.150 0.070 3.220 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.360 0.070 3.430 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.570 0.070 3.640 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.780 0.070 3.850 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.990 0.070 4.060 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.200 0.070 4.270 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.410 0.070 4.480 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.620 0.070 4.690 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.830 0.070 4.900 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.040 0.070 5.110 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.250 0.070 5.320 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.460 0.070 5.530 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.670 0.070 5.740 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.880 0.070 5.950 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.090 0.070 6.160 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.300 0.070 6.370 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.510 0.070 6.580 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.720 0.070 6.790 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.930 0.070 7.000 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.140 0.070 7.210 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.350 0.070 7.420 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.560 0.070 7.630 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.770 0.070 7.840 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.980 0.070 8.050 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.190 0.070 8.260 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.400 0.070 8.470 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.610 0.070 8.680 ;
    END
  END w_mask_in[31]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.390 0.070 12.460 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.600 0.070 12.670 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.810 0.070 12.880 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.020 0.070 13.090 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.230 0.070 13.300 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.440 0.070 13.510 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.650 0.070 13.720 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.860 0.070 13.930 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.070 0.070 14.140 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.280 0.070 14.350 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.490 0.070 14.560 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.700 0.070 14.770 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.910 0.070 14.980 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.120 0.070 15.190 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.330 0.070 15.400 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.540 0.070 15.610 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.750 0.070 15.820 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.960 0.070 16.030 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.170 0.070 16.240 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.380 0.070 16.450 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.590 0.070 16.660 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.800 0.070 16.870 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.010 0.070 17.080 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.220 0.070 17.290 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.430 0.070 17.500 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.640 0.070 17.710 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.850 0.070 17.920 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.060 0.070 18.130 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.270 0.070 18.340 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.480 0.070 18.550 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.690 0.070 18.760 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.900 0.070 18.970 ;
    END
  END rd_out[31]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.680 0.070 22.750 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.890 0.070 22.960 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.100 0.070 23.170 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.310 0.070 23.380 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.520 0.070 23.590 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.730 0.070 23.800 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.940 0.070 24.010 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.150 0.070 24.220 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.360 0.070 24.430 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.570 0.070 24.640 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.780 0.070 24.850 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.990 0.070 25.060 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.200 0.070 25.270 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.410 0.070 25.480 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.620 0.070 25.690 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.830 0.070 25.900 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.040 0.070 26.110 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.250 0.070 26.320 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.460 0.070 26.530 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.670 0.070 26.740 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.880 0.070 26.950 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.090 0.070 27.160 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.300 0.070 27.370 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.510 0.070 27.580 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.720 0.070 27.790 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.930 0.070 28.000 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.140 0.070 28.210 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.350 0.070 28.420 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.560 0.070 28.630 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.770 0.070 28.840 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.980 0.070 29.050 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.190 0.070 29.260 ;
    END
  END wd_in[31]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.970 0.070 33.040 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.180 0.070 33.250 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.390 0.070 33.460 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.600 0.070 33.670 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.810 0.070 33.880 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.020 0.070 34.090 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.230 0.070 34.300 ;
    END
  END addr_in[6]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.010 0.070 38.080 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.220 0.070 38.290 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.430 0.070 38.500 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.960 2.100 2.240 39.900 ;
      RECT 5.320 2.100 5.600 39.900 ;
      RECT 8.680 2.100 8.960 39.900 ;
      RECT 12.040 2.100 12.320 39.900 ;
      RECT 15.400 2.100 15.680 39.900 ;
      RECT 18.760 2.100 19.040 39.900 ;
      RECT 22.120 2.100 22.400 39.900 ;
      RECT 25.480 2.100 25.760 39.900 ;
      RECT 28.840 2.100 29.120 39.900 ;
      RECT 32.200 2.100 32.480 39.900 ;
      RECT 35.560 2.100 35.840 39.900 ;
      RECT 38.920 2.100 39.200 39.900 ;
      RECT 42.280 2.100 42.560 39.900 ;
      RECT 45.640 2.100 45.920 39.900 ;
      RECT 49.000 2.100 49.280 39.900 ;
      RECT 52.360 2.100 52.640 39.900 ;
      RECT 55.720 2.100 56.000 39.900 ;
      RECT 59.080 2.100 59.360 39.900 ;
      RECT 62.440 2.100 62.720 39.900 ;
      RECT 65.800 2.100 66.080 39.900 ;
      RECT 69.160 2.100 69.440 39.900 ;
      RECT 72.520 2.100 72.800 39.900 ;
      RECT 75.880 2.100 76.160 39.900 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 3.640 2.100 3.920 39.900 ;
      RECT 7.000 2.100 7.280 39.900 ;
      RECT 10.360 2.100 10.640 39.900 ;
      RECT 13.720 2.100 14.000 39.900 ;
      RECT 17.080 2.100 17.360 39.900 ;
      RECT 20.440 2.100 20.720 39.900 ;
      RECT 23.800 2.100 24.080 39.900 ;
      RECT 27.160 2.100 27.440 39.900 ;
      RECT 30.520 2.100 30.800 39.900 ;
      RECT 33.880 2.100 34.160 39.900 ;
      RECT 37.240 2.100 37.520 39.900 ;
      RECT 40.600 2.100 40.880 39.900 ;
      RECT 43.960 2.100 44.240 39.900 ;
      RECT 47.320 2.100 47.600 39.900 ;
      RECT 50.680 2.100 50.960 39.900 ;
      RECT 54.040 2.100 54.320 39.900 ;
      RECT 57.400 2.100 57.680 39.900 ;
      RECT 60.760 2.100 61.040 39.900 ;
      RECT 64.120 2.100 64.400 39.900 ;
      RECT 67.480 2.100 67.760 39.900 ;
      RECT 70.840 2.100 71.120 39.900 ;
      RECT 74.200 2.100 74.480 39.900 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 78.470 42.000 ;
    LAYER metal2 ;
    RECT 0 0 78.470 42.000 ;
    LAYER metal3 ;
    RECT 0.070 0 78.470 42.000 ;
    RECT 0 0.000 0.070 2.100 ;
    RECT 0 2.170 0.070 2.310 ;
    RECT 0 2.380 0.070 2.520 ;
    RECT 0 2.590 0.070 2.730 ;
    RECT 0 2.800 0.070 2.940 ;
    RECT 0 3.010 0.070 3.150 ;
    RECT 0 3.220 0.070 3.360 ;
    RECT 0 3.430 0.070 3.570 ;
    RECT 0 3.640 0.070 3.780 ;
    RECT 0 3.850 0.070 3.990 ;
    RECT 0 4.060 0.070 4.200 ;
    RECT 0 4.270 0.070 4.410 ;
    RECT 0 4.480 0.070 4.620 ;
    RECT 0 4.690 0.070 4.830 ;
    RECT 0 4.900 0.070 5.040 ;
    RECT 0 5.110 0.070 5.250 ;
    RECT 0 5.320 0.070 5.460 ;
    RECT 0 5.530 0.070 5.670 ;
    RECT 0 5.740 0.070 5.880 ;
    RECT 0 5.950 0.070 6.090 ;
    RECT 0 6.160 0.070 6.300 ;
    RECT 0 6.370 0.070 6.510 ;
    RECT 0 6.580 0.070 6.720 ;
    RECT 0 6.790 0.070 6.930 ;
    RECT 0 7.000 0.070 7.140 ;
    RECT 0 7.210 0.070 7.350 ;
    RECT 0 7.420 0.070 7.560 ;
    RECT 0 7.630 0.070 7.770 ;
    RECT 0 7.840 0.070 7.980 ;
    RECT 0 8.050 0.070 8.190 ;
    RECT 0 8.260 0.070 8.400 ;
    RECT 0 8.470 0.070 8.610 ;
    RECT 0 8.680 0.070 12.390 ;
    RECT 0 12.460 0.070 12.600 ;
    RECT 0 12.670 0.070 12.810 ;
    RECT 0 12.880 0.070 13.020 ;
    RECT 0 13.090 0.070 13.230 ;
    RECT 0 13.300 0.070 13.440 ;
    RECT 0 13.510 0.070 13.650 ;
    RECT 0 13.720 0.070 13.860 ;
    RECT 0 13.930 0.070 14.070 ;
    RECT 0 14.140 0.070 14.280 ;
    RECT 0 14.350 0.070 14.490 ;
    RECT 0 14.560 0.070 14.700 ;
    RECT 0 14.770 0.070 14.910 ;
    RECT 0 14.980 0.070 15.120 ;
    RECT 0 15.190 0.070 15.330 ;
    RECT 0 15.400 0.070 15.540 ;
    RECT 0 15.610 0.070 15.750 ;
    RECT 0 15.820 0.070 15.960 ;
    RECT 0 16.030 0.070 16.170 ;
    RECT 0 16.240 0.070 16.380 ;
    RECT 0 16.450 0.070 16.590 ;
    RECT 0 16.660 0.070 16.800 ;
    RECT 0 16.870 0.070 17.010 ;
    RECT 0 17.080 0.070 17.220 ;
    RECT 0 17.290 0.070 17.430 ;
    RECT 0 17.500 0.070 17.640 ;
    RECT 0 17.710 0.070 17.850 ;
    RECT 0 17.920 0.070 18.060 ;
    RECT 0 18.130 0.070 18.270 ;
    RECT 0 18.340 0.070 18.480 ;
    RECT 0 18.550 0.070 18.690 ;
    RECT 0 18.760 0.070 18.900 ;
    RECT 0 18.970 0.070 22.680 ;
    RECT 0 22.750 0.070 22.890 ;
    RECT 0 22.960 0.070 23.100 ;
    RECT 0 23.170 0.070 23.310 ;
    RECT 0 23.380 0.070 23.520 ;
    RECT 0 23.590 0.070 23.730 ;
    RECT 0 23.800 0.070 23.940 ;
    RECT 0 24.010 0.070 24.150 ;
    RECT 0 24.220 0.070 24.360 ;
    RECT 0 24.430 0.070 24.570 ;
    RECT 0 24.640 0.070 24.780 ;
    RECT 0 24.850 0.070 24.990 ;
    RECT 0 25.060 0.070 25.200 ;
    RECT 0 25.270 0.070 25.410 ;
    RECT 0 25.480 0.070 25.620 ;
    RECT 0 25.690 0.070 25.830 ;
    RECT 0 25.900 0.070 26.040 ;
    RECT 0 26.110 0.070 26.250 ;
    RECT 0 26.320 0.070 26.460 ;
    RECT 0 26.530 0.070 26.670 ;
    RECT 0 26.740 0.070 26.880 ;
    RECT 0 26.950 0.070 27.090 ;
    RECT 0 27.160 0.070 27.300 ;
    RECT 0 27.370 0.070 27.510 ;
    RECT 0 27.580 0.070 27.720 ;
    RECT 0 27.790 0.070 27.930 ;
    RECT 0 28.000 0.070 28.140 ;
    RECT 0 28.210 0.070 28.350 ;
    RECT 0 28.420 0.070 28.560 ;
    RECT 0 28.630 0.070 28.770 ;
    RECT 0 28.840 0.070 28.980 ;
    RECT 0 29.050 0.070 29.190 ;
    RECT 0 29.260 0.070 32.970 ;
    RECT 0 33.040 0.070 33.180 ;
    RECT 0 33.250 0.070 33.390 ;
    RECT 0 33.460 0.070 33.600 ;
    RECT 0 33.670 0.070 33.810 ;
    RECT 0 33.880 0.070 34.020 ;
    RECT 0 34.090 0.070 34.230 ;
    RECT 0 34.300 0.070 38.010 ;
    RECT 0 38.080 0.070 38.220 ;
    RECT 0 38.290 0.070 38.430 ;
    RECT 0 38.500 0.070 42.000 ;
    LAYER metal4 ;
    RECT 0 0 78.470 2.100 ;
    RECT 0 39.900 78.470 42.000 ;
    RECT 0.000 2.100 1.960 39.900 ;
    RECT 2.240 2.100 3.640 39.900 ;
    RECT 3.920 2.100 5.320 39.900 ;
    RECT 5.600 2.100 7.000 39.900 ;
    RECT 7.280 2.100 8.680 39.900 ;
    RECT 8.960 2.100 10.360 39.900 ;
    RECT 10.640 2.100 12.040 39.900 ;
    RECT 12.320 2.100 13.720 39.900 ;
    RECT 14.000 2.100 15.400 39.900 ;
    RECT 15.680 2.100 17.080 39.900 ;
    RECT 17.360 2.100 18.760 39.900 ;
    RECT 19.040 2.100 20.440 39.900 ;
    RECT 20.720 2.100 22.120 39.900 ;
    RECT 22.400 2.100 23.800 39.900 ;
    RECT 24.080 2.100 25.480 39.900 ;
    RECT 25.760 2.100 27.160 39.900 ;
    RECT 27.440 2.100 28.840 39.900 ;
    RECT 29.120 2.100 30.520 39.900 ;
    RECT 30.800 2.100 32.200 39.900 ;
    RECT 32.480 2.100 33.880 39.900 ;
    RECT 34.160 2.100 35.560 39.900 ;
    RECT 35.840 2.100 37.240 39.900 ;
    RECT 37.520 2.100 38.920 39.900 ;
    RECT 39.200 2.100 40.600 39.900 ;
    RECT 40.880 2.100 42.280 39.900 ;
    RECT 42.560 2.100 43.960 39.900 ;
    RECT 44.240 2.100 45.640 39.900 ;
    RECT 45.920 2.100 47.320 39.900 ;
    RECT 47.600 2.100 49.000 39.900 ;
    RECT 49.280 2.100 50.680 39.900 ;
    RECT 50.960 2.100 52.360 39.900 ;
    RECT 52.640 2.100 54.040 39.900 ;
    RECT 54.320 2.100 55.720 39.900 ;
    RECT 56.000 2.100 57.400 39.900 ;
    RECT 57.680 2.100 59.080 39.900 ;
    RECT 59.360 2.100 60.760 39.900 ;
    RECT 61.040 2.100 62.440 39.900 ;
    RECT 62.720 2.100 64.120 39.900 ;
    RECT 64.400 2.100 65.800 39.900 ;
    RECT 66.080 2.100 67.480 39.900 ;
    RECT 67.760 2.100 69.160 39.900 ;
    RECT 69.440 2.100 70.840 39.900 ;
    RECT 71.120 2.100 72.520 39.900 ;
    RECT 72.800 2.100 74.200 39.900 ;
    RECT 74.480 2.100 75.880 39.900 ;
    RECT 76.160 2.100 78.470 39.900 ;
    LAYER OVERLAP ;
    RECT 0 0 78.470 42.000 ;
  END
END fakeram45_128x32

END LIBRARY
