// //#############################################################################
// //# Function: Or-And (oa31) Gate                                              #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_oa31 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a0,
//     input  a1,
//     input  a2,
//     input  b0,
//     output z
// );
// 
//     assign z = (a0 | a1 | a2) & b0;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_oa31.v:10.1-22.10" *)
module la_oa31 (
    a0,
    a1,
    a2,
    b0,
    z
);
  wire _0_;
  (* src = "inputs/la_oa31.v:13.12-13.14" *)
  input a0;
  wire a0;
  (* src = "inputs/la_oa31.v:14.12-14.14" *)
  input a1;
  wire a1;
  (* src = "inputs/la_oa31.v:15.12-15.14" *)
  input a2;
  wire a2;
  (* src = "inputs/la_oa31.v:16.12-16.14" *)
  input b0;
  wire b0;
  (* src = "inputs/la_oa31.v:17.12-17.13" *)
  output z;
  wire z;
  sky130_fd_sc_hdll__o31ai_2 _1_ (
      .A1(a1),
      .A2(a0),
      .A3(a2),
      .B1(b0),
      .Y (_0_)
  );
  sky130_fd_sc_hdll__inv_1 _2_ (
      .A(_0_),
      .Y(z)
  );
endmodule
