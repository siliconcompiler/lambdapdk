// //#############################################################################
// //# Function:  Positive edge-triggered static inverting D-type flop-flop with #
// //             async active low reset and scan input                          #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_sdffrqn #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      si,
//     input      se,
//     input      clk,
//     input      nreset,
//     output reg qn
// );
// 
//     always @(posedge clk or negedge nreset)
//         if (!nreset) qn <= 1'b1;
//         else qn <= se ? ~si : ~d;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
module la_sdffrqn (
    d,
    si,
    se,
    clk,
    nreset,
    qn
);
  wire _0_;
  (* unused_bits = "0" *)
  wire _1_;
  (* src = "generated" *)
  input clk;
  wire clk;
  (* src = "generated" *)
  input d;
  wire d;
  (* src = "generated" *)
  input nreset;
  wire nreset;
  (* src = "generated" *)
  output qn;
  wire qn;
  (* src = "generated" *)
  input se;
  wire se;
  (* src = "generated" *)
  input si;
  wire si;
  sg13g2_mux2_1 _2_ (
      .A0(d),
      .A1(si),
      .S (se),
      .X (_0_)
  );
  (* src = "generated" *)
  sg13g2_dfrbp_1 _3_ (
      .CLK(clk),
      .D(_0_),
      .Q(_1_),
      .Q_N(qn),
      .RESET_B(nreset)
  );
endmodule
