// //#############################################################################
// //# Function: Dual data rate input buffer                                     #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_iddr #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      clk,      // clock
//     input      in,       // data input sampled on both edges of clock
//     output reg outrise,  // rising edge sample
//     output reg outfall   // falling edge sample
// );
// 
//   // Negedge Sample
//   always @(negedge clk) outfall <= in;
// 
//   // Posedge Sample
//   reg inrise;
//   always @(posedge clk) inrise <= in;
// 
//   // Posedge Latch (for hold)
//   always @(clk or inrise) if (~clk) outrise <= inrise;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_iddr.v:10.1-29.10" *)
module la_iddr (
    clk,
    in,
    outrise,
    outfall
);
  wire _0_;
  (* unused_bits = "0" *)
  wire _1_;
  (* unused_bits = "0" *)
  wire _2_;
  (* src = "inputs/la_iddr.v:13.16-13.19" *)
  input clk;
  wire clk;
  (* src = "inputs/la_iddr.v:14.16-14.18" *)
  input in;
  wire in;
  (* src = "inputs/la_iddr.v:23.7-23.13" *)
  wire inrise;
  (* src = "inputs/la_iddr.v:16.16-16.23" *)
  output outfall;
  wire outfall;
  (* src = "inputs/la_iddr.v:15.16-15.23" *)
  output outrise;
  wire outrise;
  INV_X2 _3_ (
      .A (clk),
      .ZN(_0_)
  );
  (* module_not_derived = 32'b00000000000000000000000000000001 *)
      (* src = "inputs/la_iddr.v:27.3-27.55|/home/pgadfort/lambdapdk/lambdapdk/freepdk45/libs/nangate45/techmap/yosys/cells_latch.v:13.12-17.10" *)
  DLL_X1 _4_ (
      .D (inrise),
      .GN(clk),
      .Q (outrise)
  );
  (* src = "inputs/la_iddr.v:24.3-24.38" *)
  DFF_X1 _5_ (
      .CK(clk),
      .D (in),
      .Q (inrise),
      .QN(_2_)
  );
  (* src = "inputs/la_iddr.v:20.3-20.39" *)
  DFF_X1 _6_ (
      .CK(_0_),
      .D (in),
      .Q (outfall),
      .QN(_1_)
  );
endmodule
