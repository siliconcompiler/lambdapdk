// //#############################################################################
// //# Function: Carry Save Adder (4:2) (aka 5:3)                                #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_csa42 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     input  b,
//     input  c,
//     input  d,
//     input  cin,
//     output sum,
//     output carry,
//     output cout
// );
// 
//     assign cout   = (a & b) | (b & c) | (a & c);
//     assign sumint = a ^ b ^ c;
//     assign sum    = cin ^ d ^ sumint;
//     assign carry  = (cin & d) | (cin & sumint) | (d & sumint);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
(* keep_hierarchy *)
module la_csa42 (
    a,
    b,
    c,
    d,
    cin,
    sum,
    carry,
    cout
);
  (* force_downto = 32'b00000000000000000000000000000001 *) (* src = "generated" *)
  wire _00_;
  (* force_downto = 32'b00000000000000000000000000000001 *) (* src = "generated" *)
  wire _01_;
  (* force_downto = 32'b00000000000000000000000000000001 *) (* src = "generated" *)
  wire _02_;
  (* force_downto = 32'b00000000000000000000000000000001 *) (* src = "generated" *)
  wire _03_;
  (* force_downto = 32'b00000000000000000000000000000001 *) (* src = "generated" *)
  wire _04_;
  (* force_downto = 32'b00000000000000000000000000000001 *) (* src = "generated" *)
  wire _05_;
  (* src = "generated" *)
  input a;
  wire a;
  (* src = "generated" *)
  input b;
  wire b;
  (* src = "generated" *)
  input c;
  wire c;
  (* src = "generated" *)
  output carry;
  wire carry;
  (* src = "generated" *)
  input cin;
  wire cin;
  (* src = "generated" *)
  output cout;
  wire cout;
  (* src = "generated" *)
  input d;
  wire d;
  (* src = "generated" *)
  output sum;
  wire sum;
  INVx2_ASAP7_75t_L _06_ (
      .A(a),
      .Y(_00_)
  );
  INVx2_ASAP7_75t_L _07_ (
      .A(d),
      .Y(_03_)
  );
  INVx2_ASAP7_75t_L _08_ (
      .A(b),
      .Y(_01_)
  );
  INVx2_ASAP7_75t_L _09_ (
      .A(cin),
      .Y(_04_)
  );
  INVx2_ASAP7_75t_L _10_ (
      .A(c),
      .Y(_02_)
  );
  (* module_not_derived = 32'b00000000000000000000000000000001 *) (* src = "generated" *)
  FAx1_ASAP7_75t_L _11_ (
      .A  (_00_),
      .B  (_01_),
      .CI (_02_),
      .CON(cout),
      .SN (_05_)
  );
  (* module_not_derived = 32'b00000000000000000000000000000001 *) (* src = "generated" *)
  FAx1_ASAP7_75t_L _12_ (
      .A  (_03_),
      .B  (_04_),
      .CI (_05_),
      .CON(carry),
      .SN (sum)
  );
endmodule
