// //#############################################################################
// //# Function: Positive edge-triggered static D-type flop-flop                 #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_dffq #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      clk,
//     output reg q
// );
// 
//   always @(posedge clk) q <= d;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_dffq.v:10.1-20.10" *)
module la_dffq (
    d,
    clk,
    q
);
  wire _0_;
  (* src = "inputs/la_dffq.v:14.16-14.19" *)
  input clk;
  wire clk;
  (* src = "inputs/la_dffq.v:13.16-13.17" *)
  input d;
  wire d;
  (* src = "inputs/la_dffq.v:15.16-15.17" *)
  output q;
  wire q;
  INVx2_ASAP7_75t_R _1_ (
      .A(_0_),
      .Y(q)
  );
  (* src = "inputs/la_dffq.v:18.3-18.32" *)
  DFFHQNx1_ASAP7_75t_R _2_ (
      .CLK(clk),
      .D  (d),
      .QN (_0_)
  );
endmodule
