// //#############################################################################
// //# Function:  Positive edge-triggered static inverting D-type flop-flop with #
// //             async active low set and scan input                            #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_sdffsqn #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      si,
//     input      se,
//     input      clk,
//     input      nset,
//     output reg qn
// );
// 
//     always @(posedge clk or negedge nset)
//         if (!nset) qn <= 1'b0;
//         else qn <= se ? ~si : ~d;
// 
// endmodule

/* Generated by Yosys 0.40 (git sha1 a1bb0255d, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_sdffsqn(d, si, se, clk, nset, qn);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  input clk;
  wire clk;
  input d;
  wire d;
  input nset;
  wire nset;
  output qn;
  wire qn;
  input se;
  wire se;
  input si;
  wire si;
  INVx1_ASAP7_75t_R _05_ (
    .A(si),
    .Y(_02_)
  );
  NOR2x1_ASAP7_75t_R _06_ (
    .A(d),
    .B(se),
    .Y(_03_)
  );
  AO21x1_ASAP7_75t_R _07_ (
    .A1(_02_),
    .A2(se),
    .B(_03_),
    .Y(_00_)
  );
  INVx1_ASAP7_75t_R _08_ (
    .A(_01_),
    .Y(qn)
  );
  DFFASRHQNx1_ASAP7_75t_R _09_ (
    .CLK(clk),
    .D(_00_),
    .QN(_01_),
    .RESETN(_04_),
    .SETN(nset)
  );
  TIEHIx1_ASAP7_75t_R _10_ (
    .H(_04_)
  );
endmodule
