// //#############################################################################
// //# Function: Power isolation circuit                                         #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_isolo #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  iso,  // isolation signal
//     input  in,   // input
//     output out   // out = ~iso & in
// );
// 
//     assign out = ~iso & in;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
module la_isolo (
    iso,
    in,
    out
);
  (* src = "generated" *)
  input in;
  wire in;
  (* src = "generated" *)
  input iso;
  wire iso;
  (* src = "generated" *)
  output out;
  wire out;
  sky130_fd_sc_hd__nor2b_4 _0_ (
      .A  (iso),
      .B_N(in),
      .Y  (out)
  );
endmodule
