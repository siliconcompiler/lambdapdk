// //#############################################################################
// //# Function: 4 Input Or Gate                                                 #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_or4 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     input  b,
//     input  c,
//     input  d,
//     output z
// );
// 
//     assign z = a | b | c | d;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
(* keep_hierarchy *)
module la_or4 (
    a,
    b,
    c,
    d,
    z
);
  (* src = "generated" *)
  input a;
  wire a;
  (* src = "generated" *)
  input b;
  wire b;
  (* src = "generated" *)
  input c;
  wire c;
  (* src = "generated" *)
  input d;
  wire d;
  (* src = "generated" *)
  output z;
  wire z;
  gf180mcu_fd_sc_mcu9t5v0__or4_4 _0_ (
      .A1(b),
      .A2(a),
      .A3(c),
      .A4(d),
      .Z (z)
  );
endmodule
