// //#############################################################################
// //# Function: Power isolation circuit                                         #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_isohi
//   #(parameter PROP = "DEFAULT")
//    (
//     input  iso, // isolation signal
//     input  in, // input
//     output out  // out = iso | in
//     );
// 
//    assign out = iso | in;
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_isohi(iso, in, out);
  input in;
  wire in;
  input iso;
  wire iso;
  output out;
  wire out;
  gf180mcu_fd_sc_mcu7t5v0__or2_2 _0_ (
    .A1(in),
    .A2(iso),
    .Z(out)
  );
endmodule
