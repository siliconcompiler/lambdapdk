// //#############################################################################
// //# Function: 4 Input Nor Gate                                                #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_nor4 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     input  b,
//     input  c,
//     input  d,
//     output z
// );
// 
//     assign z = ~(a | b | c | d);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_nor4.v:10.1-22.10" *)
module la_nor4 (
    a,
    b,
    c,
    d,
    z
);
  (* src = "inputs/la_nor4.v:13.12-13.13" *)
  input a;
  wire a;
  (* src = "inputs/la_nor4.v:14.12-14.13" *)
  input b;
  wire b;
  (* src = "inputs/la_nor4.v:15.12-15.13" *)
  input c;
  wire c;
  (* src = "inputs/la_nor4.v:16.12-16.13" *)
  input d;
  wire d;
  (* src = "inputs/la_nor4.v:17.12-17.13" *)
  output z;
  wire z;
  sky130_fd_sc_hd__nor4_4 _0_ (
      .A(b),
      .B(a),
      .C(c),
      .D(d),
      .Y(z)
  );
endmodule
