// //#############################################################################
// //# Function: Positive edge-triggered inverting static D-type flop-flop       #
// //#           with scan input.                                                #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_sdffqn #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      si,
//     input      se,
//     input      clk,
//     output reg qn
// );
// 
//     always @(posedge clk) qn <= se ? ~si : ~d;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
(* keep_hierarchy *)
module la_sdffqn (
    d,
    si,
    se,
    clk,
    qn
);
  (* src = "generated" *)
  wire _0_;
  wire _1_;
  wire _2_;
  wire _3_;
  (* src = "generated" *)
  input clk;
  wire clk;
  (* src = "generated" *)
  input d;
  wire d;
  (* src = "generated" *)
  output qn;
  wire qn;
  (* src = "generated" *)
  input se;
  wire se;
  (* src = "generated" *)
  input si;
  wire si;
  INVx1_ASAP7_75t_R _4_ (
      .A(si),
      .Y(_2_)
  );
  NOR2x1_ASAP7_75t_R _5_ (
      .A(d),
      .B(se),
      .Y(_3_)
  );
  AO21x1_ASAP7_75t_R _6_ (
      .A1(_2_),
      .A2(se),
      .B (_3_),
      .Y (_0_)
  );
  INVx1_ASAP7_75t_R _7_ (
      .A(_1_),
      .Y(qn)
  );
  (* src = "generated" *)
  DFFHQNx1_ASAP7_75t_R _8_ (
      .CLK(clk),
      .D  (_0_),
      .QN (_1_)
  );
endmodule
