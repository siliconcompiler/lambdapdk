// //#############################################################################
// //# Function: 2-Input AND Gate                                                #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_and2 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     input  b,
//     output z
// );
// 
//     assign z = a & b;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
module la_and2 (
    a,
    b,
    z
);
  (* src = "generated" *)
  input a;
  wire a;
  (* src = "generated" *)
  input b;
  wire b;
  (* src = "generated" *)
  output z;
  wire z;
  AND2x4_ASAP7_75t_R _0_ (
      .A(b),
      .B(a),
      .Y(z)
  );
endmodule
