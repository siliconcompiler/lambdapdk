// //#############################################################################
// //# Function: And-Or (ao32) Gate                                              #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_ao32 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a0,
//     input  a1,
//     input  a2,
//     input  b0,
//     input  b1,
//     output z
// );
// 
//     assign z = (a0 & a1 & a2) | (b0 & b1);
// 
// endmodule

/* Generated by Yosys 0.40+33 (git sha1 cd1fb8b15, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_ao32(a0, a1, a2, b0, b1, z);
  wire _0_;
  wire _1_;
  input a0;
  wire a0;
  input a1;
  wire a1;
  input a2;
  wire a2;
  input b0;
  wire b0;
  input b1;
  wire b1;
  output z;
  wire z;
  sg13g2_nand2_1 _2_ (
    .A(b1),
    .B(b0),
    .Y(_0_)
  );
  sg13g2_nand3_1 _3_ (
    .A(a1),
    .B(a0),
    .C(a2),
    .Y(_1_)
  );
  sg13g2_nand2_1 _4_ (
    .A(_0_),
    .B(_1_),
    .Y(z)
  );
endmodule
