// //#############################################################################
// //# Function: 4-Input Inverting Mux                                           #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_muxi4 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  d0,
//     input  d1,
//     input  d2,
//     input  d3,
//     input  s0,
//     input  s1,
//     output z
// );
// 
//     assign z = ~((d0 & ~s1 & ~s0) | (d1 & ~s1 & s0) | (d2 & s1 & ~s0) | (d3 & s1 & s0));
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
module la_muxi4 (
    d0,
    d1,
    d2,
    d3,
    s0,
    s1,
    z
);
  wire _0_;
  wire _1_;
  (* src = "generated" *)
  input d0;
  wire d0;
  (* src = "generated" *)
  input d1;
  wire d1;
  (* src = "generated" *)
  input d2;
  wire d2;
  (* src = "generated" *)
  input d3;
  wire d3;
  (* src = "generated" *)
  input s0;
  wire s0;
  (* src = "generated" *)
  input s1;
  wire s1;
  (* src = "generated" *)
  output z;
  wire z;
  sky130_fd_sc_hdll__mux2i_1 _2_ (
      .A0(d0),
      .A1(d1),
      .S (s0),
      .Y (_0_)
  );
  sky130_fd_sc_hdll__mux2i_1 _3_ (
      .A0(d2),
      .A1(d3),
      .S (s0),
      .Y (_1_)
  );
  sky130_fd_sc_hdll__clkmux2_1 _4_ (
      .A0(_0_),
      .A1(_1_),
      .S (s1),
      .X (z)
  );
endmodule
