// //#############################################################################
// //# Function: Carry Save Adder (4:2) (aka 5:3)                                #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_csa42 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     input  b,
//     input  c,
//     input  d,
//     input  cin,
//     output sum,
//     output carry,
//     output cout
// );
// 
//     assign cout   = (a & b) | (b & c) | (a & c);
//     assign sumint = a ^ b ^ c;
//     assign sum    = cin ^ d ^ sumint;
//     assign carry  = (cin & d) | (cin & sumint) | (d & sumint);
// 
// endmodule

/* Generated by Yosys 0.40 (git sha1 a1bb0255d, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_csa42(a, b, c, d, cin, sum, carry, cout);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  input a;
  wire a;
  input b;
  wire b;
  input c;
  wire c;
  output carry;
  wire carry;
  input cin;
  wire cin;
  output cout;
  wire cout;
  input d;
  wire d;
  output sum;
  wire sum;
  INVx1_ASAP7_75t_L _06_ (
    .A(a),
    .Y(_00_)
  );
  INVx1_ASAP7_75t_L _07_ (
    .A(d),
    .Y(_03_)
  );
  INVx1_ASAP7_75t_L _08_ (
    .A(b),
    .Y(_01_)
  );
  INVx1_ASAP7_75t_L _09_ (
    .A(cin),
    .Y(_04_)
  );
  INVx1_ASAP7_75t_L _10_ (
    .A(c),
    .Y(_02_)
  );
  FAx1_ASAP7_75t_L _11_ (
    .A(_00_),
    .B(_01_),
    .CI(_02_),
    .CON(cout),
    .SN(_05_)
  );
  FAx1_ASAP7_75t_L _12_ (
    .A(_03_),
    .B(_04_),
    .CI(_05_),
    .CON(carry),
    .SN(sum)
  );
endmodule
