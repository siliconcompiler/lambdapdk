// //#############################################################################
// //# Function: And-Or-Inverter (aoi31) Gate                                    #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_aoi31 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a0,
//     input  a1,
//     input  a2,
//     input  b0,
//     output z
// );
// 
//     assign z = ~((a0 & a1 & a2) | b0);
// 
// endmodule

/* Generated by Yosys 0.40+33 (git sha1 cd1fb8b15, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_aoi31(a0, a1, a2, b0, z);
  wire _0_;
  input a0;
  wire a0;
  input a1;
  wire a1;
  input a2;
  wire a2;
  input b0;
  wire b0;
  output z;
  wire z;
  sg13g2_nand3_1 _1_ (
    .A(a1),
    .B(a0),
    .C(a2),
    .Y(_0_)
  );
  sg13g2_nor2b_1 _2_ (
    .A(b0),
    .B_N(_0_),
    .Y(z)
  );
endmodule
