// //#############################################################################
// //# Function: Clock Inverter                                                  #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_clkinv #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     output z
// );
// 
//     assign z = ~a;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
module la_clkinv (
    a,
    z
);
  (* src = "generated" *)
  input a;
  wire a;
  (* src = "generated" *)
  output z;
  wire z;
  INVx2_ASAP7_75t_R _0_ (
      .A(a),
      .Y(z)
  );
endmodule
