// //#############################################################################
// //# Function: Inverter                                                        #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_inv #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     output z
// );
// 
//     assign z = ~a;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_inv.v:10.1-19.10" *)
module la_inv (
    a,
    z
);
  (* src = "inputs/la_inv.v:13.12-13.13" *)
  input a;
  wire a;
  (* src = "inputs/la_inv.v:14.12-14.13" *)
  output z;
  wire z;
  sg13g2_inv_2 _0_ (
      .A(a),
      .Y(z)
  );
endmodule
