// //#############################################################################
// //# Function: Positive edge-triggered inverting static D-type flop-flop       #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_dffqn #(
//     parameter PROP = "DEFAULT"
// ) (
//     input d,
//     input clk,
//     output reg qn
// );
// 
//     always @(posedge clk) qn <= ~d;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
(* keep_hierarchy *)
module la_dffqn (
    d,
    clk,
    qn
);
  (* src = "generated" *)
  wire _0_;
  wire _1_;
  (* src = "generated" *)
  input clk;
  wire clk;
  (* src = "generated" *)
  input d;
  wire d;
  (* src = "generated" *)
  output qn;
  wire qn;
  INVx2_ASAP7_75t_L _2_ (
      .A(d),
      .Y(_0_)
  );
  INVx2_ASAP7_75t_L _3_ (
      .A(_1_),
      .Y(qn)
  );
  (* src = "generated" *)
  DFFHQNx1_ASAP7_75t_L _4_ (
      .CLK(clk),
      .D  (_0_),
      .QN (_1_)
  );
endmodule
