# Copyright 2024 ZeroASIC Corp
# 
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
# 
#      https://www.apache.org/licenses/LICENSE-2.0
# 
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER metal1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 1.6 ;
  SPACING 0.8 ;
  WIDTH 0.8 ;
  MAXWIDTH 5.0 ;
END metal1

LAYER via1
  TYPE CUT ;
  SPACING 0.4 ;
  WIDTH 0.4 ;
END via1

LAYER metal2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 1.6 ;
  SPACING 0.8 ;
  WIDTH 0.8 ;
  MAXWIDTH 5.0 ;
END metal2

LAYER via2
  TYPE CUT ;
  SPACING 0.4 ;
  WIDTH 0.4 ;
END via2

LAYER metal3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 1.6 ;
  SPACING 0.8 ;
  WIDTH 0.8 ;
  MAXWIDTH 5.0 ;
END metal3

LAYER via3
  TYPE CUT ;
  SPACING 0.4 ;
  WIDTH 0.4 ;
END via3

LAYER metal4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 1.6 ;
  SPACING 0.8 ;
  WIDTH 0.8 ;
  MAXWIDTH 5.0 ;
END metal4

LAYER via4
  TYPE CUT ;
  SPACING 0.4 ;
  WIDTH 0.4 ;
END via4

LAYER topmetal
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 1.6 ;
  SPACING 0.8 ;
  WIDTH 0.8 ;
END topmetal

VIA VIA1_1 DEFAULT
  LAYER via1 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER metal1 ;
    RECT -0.600 -0.600 0.600 0.600 ;
  LAYER metal2 ;
    RECT -0.600 -0.600 0.600 0.600 ;
END VIA1_1

VIA VIA2_1 DEFAULT
  LAYER via2 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER metal2 ;
    RECT -0.600 -0.600 0.600 0.600 ;
  LAYER metal3 ;
    RECT -0.600 -0.600 0.600 0.600 ;
END VIA2_1

VIA VIA3_1 DEFAULT
  LAYER via3 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER metal3 ;
    RECT -0.600 -0.600 0.600 0.600 ;
  LAYER metal4 ;
    RECT -0.600 -0.600 0.600 0.600 ;
END VIA3_1

VIA VIA4_1 DEFAULT
  LAYER via4 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER metal4 ;
    RECT -0.600 -0.600 0.600 0.600 ;
  LAYER topmetal ;
    RECT -0.600 -0.600 0.600 0.600 ;
END VIA4_1


SITE dummy_site
  SYMMETRY X Y ;
  CLASS core ;
  SIZE 1.0 BY 1.0 ;
END dummy_site