// //#############################################################################
// //# Function: Dual data rate input buffer                                     #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_iddr #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      clk,      // clock
//     input      in,       // data input sampled on both edges of clock
//     output reg outrise,  // rising edge sample
//     output reg outfall   // falling edge sample
// );
// 
//     // Negedge Sample
//     always @(negedge clk) outfall <= in;
// 
//     // Posedge Sample
//     reg inrise;
//     always @(posedge clk) inrise <= in;
// 
//     // Posedge Latch (for hold)
//     always @(clk or inrise) if (~clk) outrise <= inrise;
// 
// endmodule

/* Generated by Yosys 0.41 (git sha1 c1ad37779, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_iddr(clk, in, outrise, outfall);
  wire _0_;
  wire _1_;
  input clk;
  wire clk;
  input in;
  wire in;
  wire inrise;
  output outfall;
  wire outfall;
  output outrise;
  wire outrise;
  sky130_fd_sc_hdll__inv_2 _2_ (
    .A(clk),
    .Y(_0_)
  );
  sky130_fd_sc_hdll__dlxtn_1 _3_ (
    .D(inrise),
    .GATE_N(clk),
    .Q(outrise)
  );
  sky130_fd_sc_hdll__dfrtp_1 _4_ (
    .CLK(clk),
    .D(in),
    .Q(inrise),
    .RESET_B(_1_)
  );
  sky130_fd_sc_hdll__dfrtp_1 _5_ (
    .CLK(_0_),
    .D(in),
    .Q(outfall),
    .RESET_B(_1_)
  );
  sky130_fd_sc_hdll__conb_1 _6_ (
    .HI(_1_)
  );
endmodule
