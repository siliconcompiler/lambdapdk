// //#############################################################################
// //# Function: 3-Input Inverting Mux                                           #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_muxi3 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  d0,
//     input  d1,
//     input  d2,
//     input  s0,
//     input  s1,
//     output z
// );
// 
//     assign z = ~((d0 & ~s0 & ~s1) | (d1 & s0 & ~s1) | (d2 & s1));
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_muxi3.v:10.1-23.10" *)
module la_muxi3 (
    d0,
    d1,
    d2,
    s0,
    s1,
    z
);
  wire _0_;
  wire _1_;
  (* src = "inputs/la_muxi3.v:13.12-13.14" *)
  input d0;
  wire d0;
  (* src = "inputs/la_muxi3.v:14.12-14.14" *)
  input d1;
  wire d1;
  (* src = "inputs/la_muxi3.v:15.12-15.14" *)
  input d2;
  wire d2;
  (* src = "inputs/la_muxi3.v:16.12-16.14" *)
  input s0;
  wire s0;
  (* src = "inputs/la_muxi3.v:17.12-17.14" *)
  input s1;
  wire s1;
  (* src = "inputs/la_muxi3.v:18.12-18.13" *)
  output z;
  wire z;
  sg13g2_mux2_1 _2_ (
      .A0(d0),
      .A1(d1),
      .S (s0),
      .X (_0_)
  );
  sg13g2_nand2b_1 _3_ (
      .A_N(d2),
      .B  (s1),
      .Y  (_1_)
  );
  sg13g2_o21ai_1 _4_ (
      .A1(s1),
      .A2(_0_),
      .B1(_1_),
      .Y (z)
  );
endmodule
