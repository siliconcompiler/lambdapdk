// //#############################################################################
// //# Function: 3-Input one-hot mux                                             #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_dmux3 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  sel0,
//     input  sel1,
//     input  sel2,
//     input  in0,
//     input  in1,
//     input  in2,
//     output out
// );
// 
//   assign out = (sel0 & in0) | (sel1 & in1) | (sel2 & in2);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_dmux3.v:10.1-24.10" *)
module la_dmux3 (
    sel0,
    sel1,
    sel2,
    in0,
    in1,
    in2,
    out
);
  wire _0_;
  (* src = "inputs/la_dmux3.v:16.12-16.15" *)
  input in0;
  wire in0;
  (* src = "inputs/la_dmux3.v:17.12-17.15" *)
  input in1;
  wire in1;
  (* src = "inputs/la_dmux3.v:18.12-18.15" *)
  input in2;
  wire in2;
  (* src = "inputs/la_dmux3.v:19.12-19.15" *)
  output out;
  wire out;
  (* src = "inputs/la_dmux3.v:13.12-13.16" *)
  input sel0;
  wire sel0;
  (* src = "inputs/la_dmux3.v:14.12-14.16" *)
  input sel1;
  wire sel1;
  (* src = "inputs/la_dmux3.v:15.12-15.16" *)
  input sel2;
  wire sel2;
  AOI222_X2 _1_ (
      .A1(in2),
      .A2(sel2),
      .B1(in0),
      .B2(sel0),
      .C1(in1),
      .C2(sel1),
      .ZN(_0_)
  );
  INV_X1 _2_ (
      .A (_0_),
      .ZN(out)
  );
endmodule
