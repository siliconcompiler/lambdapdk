// //#############################################################################
// //# Function: Integrated "Or" Clock Gating Cell                               #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_clkicgor #(parameter PROP = "DEFAULT")  (
//    input  clk,// clock input
//    input  te, // test enable
//    input  en, // enable
//    output eclk  // enabled clock output
//    );
// 
//    reg 	  en_stable;
// 
//    always @ (clk or en or te)
//      if (clk)
//        en_stable <= en | te;
// 
//    assign eclk =  clk | ~en_stable;
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_clkicgor(clk, te, en, eclk);
  wire _0_;
  input clk;
  wire clk;
  output eclk;
  wire eclk;
  input en;
  wire en;
  wire en_stable;
  input te;
  wire te;
  sky130_fd_sc_hdll__or2_0 _1_ (
    .A(te),
    .B(en),
    .X(_0_)
  );
  sky130_fd_sc_hdll__nand2b_1 _2_ (
    .A_N(clk),
    .B(en_stable),
    .Y(eclk)
  );
  sky130_fd_sc_hdll__dlxtp_1 _3_ (
    .D(_0_),
    .GATE(clk),
    .Q(en_stable)
  );
endmodule
