// //#############################################################################
// //# Function: Or-And-Inverter (oai222) Gate                                   #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_oai222 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a0,
//     input  a1,
//     input  b0,
//     input  b1,
//     input  c0,
//     input  c1,
//     output z
// );
// 
//     assign z = ~((a0 | a1) & (b0 | b1) & (c0 | c1));
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
(* keep_hierarchy *)
module la_oai222 (
    a0,
    a1,
    b0,
    b1,
    c0,
    c1,
    z
);
  wire _0_;
  (* src = "generated" *)
  input a0;
  wire a0;
  (* src = "generated" *)
  input a1;
  wire a1;
  (* src = "generated" *)
  input b0;
  wire b0;
  (* src = "generated" *)
  input b1;
  wire b1;
  (* src = "generated" *)
  input c0;
  wire c0;
  (* src = "generated" *)
  input c1;
  wire c1;
  (* src = "generated" *)
  output z;
  wire z;
  sky130_fd_sc_hd__o22a_1 _1_ (
      .A1(c1),
      .A2(c0),
      .B1(a1),
      .B2(a0),
      .X (_0_)
  );
  sky130_fd_sc_hd__o21ai_2 _2_ (
      .A1(b1),
      .A2(b0),
      .B1(_0_),
      .Y (z)
  );
endmodule
