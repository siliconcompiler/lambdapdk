// //#############################################################################
// //# Function: 4-Input one-hot mux                                             #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_dmux4 #(
//     parameter PROP = "DEFAULT"  // cell property
// ) (
//     input  sel3,
//     input  sel2,
//     input  sel1,
//     input  sel0,
//     input  in3,
//     input  in2,
//     input  in1,
//     input  in0,
//     output out
// );
// 
//     assign out = (sel0 & in0) | (sel1 & in1) | (sel2 & in2) | (sel3 & in3);
// 
// endmodule

/* Generated by Yosys 0.38+92 (git sha1 84116c9a3, x86_64-conda-linux-gnu-cc 11.2.0 -fvisibility-inlines-hidden -fmessage-length=0 -march=nocona -mtune=haswell -ftree-vectorize -fPIC -fstack-protector-strong -fno-plt -O2 -ffunction-sections -fdebug-prefix-map=/root/conda-eda/conda-eda/workdir/conda-env/conda-bld/yosys_1708682838165/work=/usr/local/src/conda/yosys-0.38_93_g84116c9a3 -fdebug-prefix-map=/user/projekt_pia/miniconda3/envs/sc=/usr/local/src/conda-prefix -fPIC -Os -fno-merge-constants) */

module la_dmux4(sel3, sel2, sel1, sel0, in3, in2, in1, in0, out);
  wire _0_;
  wire _1_;
  input in0;
  wire in0;
  input in1;
  wire in1;
  input in2;
  wire in2;
  input in3;
  wire in3;
  output out;
  wire out;
  input sel0;
  wire sel0;
  input sel1;
  wire sel1;
  input sel2;
  wire sel2;
  input sel3;
  wire sel3;
  sky130_fd_sc_hdll__a22oi_2 _2_ (
    .A1(in0),
    .A2(sel0),
    .B1(in2),
    .B2(sel2),
    .Y(_0_)
  );
  sky130_fd_sc_hdll__a22oi_2 _3_ (
    .A1(in1),
    .A2(sel1),
    .B1(in3),
    .B2(sel3),
    .Y(_1_)
  );
  sky130_fd_sc_hdll__nand2_1 _4_ (
    .A(_0_),
    .B(_1_),
    .Y(out)
  );
endmodule
