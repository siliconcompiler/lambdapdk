// //#############################################################################
// //# Function: Carry Save Adder (3:2)                                          #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_csa32 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     input  b,
//     input  c,
//     output sum,
//     output carry
// );
// 
//     assign sum   = a ^ b ^ c;
//     assign carry = (a & b) | (b & c) | (c & a);
// 
// endmodule

/* Generated by Yosys 0.38+92 (git sha1 84116c9a3, x86_64-conda-linux-gnu-cc 11.2.0 -fvisibility-inlines-hidden -fmessage-length=0 -march=nocona -mtune=haswell -ftree-vectorize -fPIC -fstack-protector-strong -fno-plt -O2 -ffunction-sections -fdebug-prefix-map=/root/conda-eda/conda-eda/workdir/conda-env/conda-bld/yosys_1708682838165/work=/usr/local/src/conda/yosys-0.38_93_g84116c9a3 -fdebug-prefix-map=/user/projekt_pia/miniconda3/envs/sc=/usr/local/src/conda-prefix -fPIC -Os -fno-merge-constants) */

module la_csa32(a, b, c, sum, carry);
  wire _0_;
  wire _1_;
  wire _2_;
  input a;
  wire a;
  input b;
  wire b;
  input c;
  wire c;
  output carry;
  wire carry;
  output sum;
  wire sum;
  sky130_fd_sc_hdll__xnor2_2 _3_ (
    .A(b),
    .B(c),
    .Y(_0_)
  );
  sky130_fd_sc_hdll__xnor2_1 _4_ (
    .A(a),
    .B(_0_),
    .Y(sum)
  );
  sky130_fd_sc_hdll__nand2_1 _5_ (
    .A(b),
    .B(c),
    .Y(_1_)
  );
  sky130_fd_sc_hdll__o21ai_1 _6_ (
    .A1(b),
    .A2(c),
    .B1(a),
    .Y(_2_)
  );
  sky130_fd_sc_hdll__nand2_1 _7_ (
    .A(_1_),
    .B(_2_),
    .Y(carry)
  );
endmodule
