// //#############################################################################
// //# Function: Positive edge-triggered static D-type flop-flop with scan input #
// //#                                                                           #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_sdffq #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      si,
//     input      se,
//     input      clk,
//     output reg q
// );
// 
//     always @(posedge clk) q <= se ? si : d;
// 
// endmodule

/* Generated by Yosys 0.40 (git sha1 a1bb0255d, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_sdffq(d, si, se, clk, q);
  wire _0_;
  wire _1_;
  wire _2_;
  wire _3_;
  input clk;
  wire clk;
  input d;
  wire d;
  output q;
  wire q;
  input se;
  wire se;
  input si;
  wire si;
  INVx1_ASAP7_75t_R _4_ (
    .A(se),
    .Y(_2_)
  );
  AND2x4_ASAP7_75t_R _5_ (
    .A(si),
    .B(se),
    .Y(_3_)
  );
  AO21x1_ASAP7_75t_R _6_ (
    .A1(d),
    .A2(_2_),
    .B(_3_),
    .Y(_0_)
  );
  INVx1_ASAP7_75t_R _7_ (
    .A(_1_),
    .Y(q)
  );
  DFFHQNx1_ASAP7_75t_R _8_ (
    .CLK(clk),
    .D(_0_),
    .QN(_1_)
  );
endmodule
