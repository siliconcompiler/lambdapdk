// //#############################################################################
// //# Function: Integrated "And" Clock Gating Cell (And)                        #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_clkicgand #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  clk,  // clock input
//     input  te,   // test enable
//     input  en,   // enable (from positive edge FF)
//     output eclk  // enabled clock output
// );
// 
//     reg en_stable;
// 
//     always @(clk or en or te) if (~clk) en_stable <= en | te;
// 
//     assign eclk = clk & en_stable;
// 
// endmodule

/* Generated by Yosys 0.40 (git sha1 a1bb0255d, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_clkicgand(clk, te, en, eclk);
  wire _0_;
  input clk;
  wire clk;
  output eclk;
  wire eclk;
  input en;
  wire en;
  wire en_stable;
  input te;
  wire te;
  AND2x2_ASAP7_75t_L _1_ (
    .A(en_stable),
    .B(clk),
    .Y(eclk)
  );
  OR2x2_ASAP7_75t_L _2_ (
    .A(te),
    .B(en),
    .Y(_0_)
  );
  DLLx1_ASAP7_75t_L _3_ (
    .CLK(clk),
    .D(_0_),
    .Q(en_stable)
  );
endmodule
