// //#############################################################################
// //# Function: Negative edge-triggered static D-type flop-flop                 #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_dffnq #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      clk,
//     output reg q
// );
// 
//   always @(negedge clk) q <= d;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_dffnq.v:10.1-20.10" *)
module la_dffnq (
    d,
    clk,
    q
);
  wire _0_;
  (* src = "inputs/la_dffnq.v:14.16-14.19" *)
  input clk;
  wire clk;
  (* src = "inputs/la_dffnq.v:13.16-13.17" *)
  input d;
  wire d;
  (* src = "inputs/la_dffnq.v:15.16-15.17" *)
  output q;
  wire q;
  INVx2_ASAP7_75t_L _1_ (
      .A(_0_),
      .Y(q)
  );
  (* src = "inputs/la_dffnq.v:18.3-18.32" *)
  DFFLQNx1_ASAP7_75t_L _2_ (
      .CLK(clk),
      .D  (d),
      .QN (_0_)
  );
endmodule
