// //#############################################################################
// //# Function: Synchronizer                                                    #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_dsync #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  clk,  // clock
//     input  in,   // input data
//     output out   // synchronized data
// );
// 
//     localparam STAGES = 2;
//     localparam RND = 1;
// 
//     reg     [STAGES:0] shiftreg;
//     integer            sync_delay;
// 
//     always @(posedge clk) begin
//         shiftreg[STAGES:0] <= {shiftreg[STAGES-1:0], in};
// `ifndef SYNTHESIS
//         sync_delay <= {$random} % 2;
// `endif
//     end
// 
// `ifdef SYNTHESIS
//     assign out = shiftreg[STAGES-1];
// `else
//     assign out = (|sync_delay & (|RND)) ? shiftreg[STAGES] : shiftreg[STAGES-1];
// `endif
// 
// endmodule

/* Generated by Yosys 0.40 (git sha1 a1bb0255d, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_dsync(clk, in, out);
  wire _0_;
  wire _1_;
  input clk;
  wire clk;
  input in;
  wire in;
  output out;
  wire out;
  wire \shiftreg[0] ;
  INVx1_ASAP7_75t_SL _2_ (
    .A(_0_),
    .Y(out)
  );
  INVx1_ASAP7_75t_SL _3_ (
    .A(_1_),
    .Y(\shiftreg[0] )
  );
  DFFHQNx1_ASAP7_75t_SL _4_ (
    .CLK(clk),
    .D(in),
    .QN(_1_)
  );
  DFFHQNx1_ASAP7_75t_SL _5_ (
    .CLK(clk),
    .D(\shiftreg[0] ),
    .QN(_0_)
  );
endmodule
