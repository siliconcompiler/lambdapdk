// //#############################################################################
// //# Function:  Positive edge-triggered static inverting D-type flop-flop with #
// //             async active low reset and scan input                          #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_sdffrqn #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      si,
//     input      se,
//     input      clk,
//     input      nreset,
//     output reg qn
// );
// 
//     always @(posedge clk or negedge nreset)
//         if (!nreset) qn <= 1'b1;
//         else qn <= se ? ~si : ~d;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_sdffrqn.v:11.1-26.10" *)
module la_sdffrqn (
    d,
    si,
    se,
    clk,
    nreset,
    qn
);
  wire _0_;
  (* unused_bits = "0" *)
  wire _1_;
  (* src = "inputs/la_sdffrqn.v:17.16-17.19" *)
  input clk;
  wire clk;
  (* src = "inputs/la_sdffrqn.v:14.16-14.17" *)
  input d;
  wire d;
  (* src = "inputs/la_sdffrqn.v:18.16-18.22" *)
  input nreset;
  wire nreset;
  (* src = "inputs/la_sdffrqn.v:19.16-19.18" *)
  output qn;
  wire qn;
  (* src = "inputs/la_sdffrqn.v:16.16-16.18" *)
  input se;
  wire se;
  (* src = "inputs/la_sdffrqn.v:15.16-15.18" *)
  input si;
  wire si;
  sg13g2_mux2_1 _2_ (
      .A0(d),
      .A1(si),
      .S (se),
      .X (_0_)
  );
  (* src = "inputs/la_sdffrqn.v:22.5-24.34" *)
  sg13g2_dfrbp_1 _3_ (
      .CLK(clk),
      .D(_0_),
      .Q(_1_),
      .Q_N(qn),
      .RESET_B(nreset)
  );
endmodule
