// //#############################################################################
// //# Function:  D-type active-high transparent latch                           #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_latq #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      clk,
//     output reg q
// );
// 
//   always @(clk or d) if (clk) q <= d;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_latq.v:10.1-20.10" *)
module la_latq (
    d,
    clk,
    q
);
  (* src = "inputs/la_latq.v:14.16-14.19" *)
  input clk;
  wire clk;
  (* src = "inputs/la_latq.v:13.16-13.17" *)
  input d;
  wire d;
  (* src = "inputs/la_latq.v:15.16-15.17" *)
  output q;
  wire q;
  (* module_not_derived = 32'b00000000000000000000000000000001 *)
      (* src = "inputs/la_latq.v:18.3-18.38|/home/pgadfort/lambdapdk/lambdapdk/gf180/libs/gf180mcu_fd_sc_mcu7t5v0/techmap/yosys/cells_latch.v:2.37-6.10" *)
  gf180mcu_fd_sc_mcu7t5v0__latq_1 _0_ (
      .D(d),
      .E(clk),
      .Q(q)
  );
endmodule
