// //#############################################################################
// //# Function: Non-inverting Delay Cell                                        #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_delay #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     output z
// );
// 
//     assign z = a;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_delay.v:10.1-19.10" *)
module la_delay (
    a,
    z
);
  (* src = "inputs/la_delay.v:13.12-13.13" *)
  input a;
  wire a;
  (* src = "inputs/la_delay.v:14.12-14.13" *)
  output z;
  wire z;
  assign z = a;
endmodule
