// //#############################################################################
// //# Function: And-Or-Inverter (aoi32) Gate                                    #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_aoi32 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a0,
//     input  a1,
//     input  a2,
//     input  b0,
//     input  b1,
//     output z
// );
// 
//   assign z = ~((a0 & a1 & a2) | (b0 & b1));
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_aoi32.v:10.1-23.10" *)
module la_aoi32 (
    a0,
    a1,
    a2,
    b0,
    b1,
    z
);
  wire _0_;
  (* src = "inputs/la_aoi32.v:13.12-13.14" *)
  input a0;
  wire a0;
  (* src = "inputs/la_aoi32.v:14.12-14.14" *)
  input a1;
  wire a1;
  (* src = "inputs/la_aoi32.v:15.12-15.14" *)
  input a2;
  wire a2;
  (* src = "inputs/la_aoi32.v:16.12-16.14" *)
  input b0;
  wire b0;
  (* src = "inputs/la_aoi32.v:17.12-17.14" *)
  input b1;
  wire b1;
  (* src = "inputs/la_aoi32.v:18.12-18.13" *)
  output z;
  wire z;
  AO32x1_ASAP7_75t_SL _1_ (
      .A1(a1),
      .A2(a0),
      .A3(a2),
      .B1(b1),
      .B2(b0),
      .Y (_0_)
  );
  INVx2_ASAP7_75t_SL _2_ (
      .A(_0_),
      .Y(z)
  );
endmodule
