// //#############################################################################
// //# Function: 3-Input Mux                                                     #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_mux3 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  d0,
//     input  d1,
//     input  d2,
//     input  s0,
//     input  s1,
//     output z
// );
// 
//     assign z = (d0 & ~s0 & ~s1) | (d1 & s0 & ~s1) | (d2 & s1);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
module la_mux3 (
    d0,
    d1,
    d2,
    s0,
    s1,
    z
);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  (* src = "generated" *)
  input d0;
  wire d0;
  (* src = "generated" *)
  input d1;
  wire d1;
  (* src = "generated" *)
  input d2;
  wire d2;
  (* src = "generated" *)
  input s0;
  wire s0;
  (* src = "generated" *)
  input s1;
  wire s1;
  (* src = "generated" *)
  output z;
  wire z;
  INVx1_ASAP7_75t_L _05_ (
      .A(s1),
      .Y(_02_)
  );
  INVx1_ASAP7_75t_L _06_ (
      .A(s0),
      .Y(_03_)
  );
  AND2x2_ASAP7_75t_L _07_ (
      .A(s0),
      .B(d1),
      .Y(_04_)
  );
  AO21x1_ASAP7_75t_L _08_ (
      .A1(_03_),
      .A2(d0),
      .B (_04_),
      .Y (_00_)
  );
  AND2x2_ASAP7_75t_L _09_ (
      .A(s1),
      .B(d2),
      .Y(_01_)
  );
  AO21x1_ASAP7_75t_L _10_ (
      .A1(_02_),
      .A2(_00_),
      .B (_01_),
      .Y (z)
  );
endmodule
