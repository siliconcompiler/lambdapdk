// //#############################################################################
// //# Function: Positive edge-triggered static D-type flop-flop with scan input #
// //#                                                                           #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_sdffq #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      si,
//     input      se,
//     input      clk,
//     output reg q
// );
// 
//     always @(posedge clk) q <= se ? si : d;
// 
// endmodule

/* Generated by Yosys 0.40+33 (git sha1 cd1fb8b15, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_sdffq(d, si, se, clk, q);
  wire _0_;
  wire _1_;
  wire _2_;
  input clk;
  wire clk;
  input d;
  wire d;
  output q;
  wire q;
  input se;
  wire se;
  input si;
  wire si;
  sg13g2_mux2_1 _3_ (
    .A0(d),
    .A1(si),
    .S(se),
    .X(_0_)
  );
  sg13g2_dfrbp_1 _4_ (
    .CLK(clk),
    .D(_0_),
    .Q(q),
    .Q_N(_1_),
    .RESET_B(_2_)
  );
  sg13g2_tiehi _5_ (
    .L_HI(_2_)
  );
endmodule
