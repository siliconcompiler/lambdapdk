// //#############################################################################
// //# Function: Dual data rate output buffer                                    #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_oddr #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  clk,  // clock input
//     input  in0,  // data for clk=0
//     input  in1,  // data for clk=1
//     output out   // dual data rate output
// );
// 
//   //Making in1 stable for clk=1
//   reg in1_sh;
//   always @(clk or in1) if (~clk) in1_sh <= in1;
// 
//   //Using clock as data selector
//   assign out = clk ? in1_sh : in0;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_oddr.v:10.1-26.10" *)
module la_oddr (
    clk,
    in0,
    in1,
    out
);
  (* src = "inputs/la_oddr.v:13.12-13.15" *)
  input clk;
  wire clk;
  (* src = "inputs/la_oddr.v:14.12-14.15" *)
  input in0;
  wire in0;
  (* src = "inputs/la_oddr.v:15.12-15.15" *)
  input in1;
  wire in1;
  (* src = "inputs/la_oddr.v:20.7-20.13" *)
  wire in1_sh;
  (* src = "inputs/la_oddr.v:16.12-16.15" *)
  output out;
  wire out;
  sky130_fd_sc_hdll__clkmux2_1 _0_ (
      .A0(in0),
      .A1(in1_sh),
      .S (clk),
      .X (out)
  );
  (* module_not_derived = 32'b00000000000000000000000000000001 *)
      (* src = "inputs/la_oddr.v:21.3-21.48|/home/pgadfort/lambdapdk/lambdapdk/sky130/libs/sky130hdll/techmap/yosys/cells_latch.v:2.32-6.10" *)
  sky130_fd_sc_hdll__dlxtn_1 _1_ (
      .D(in1),
      .GATE_N(clk),
      .Q(in1_sh)
  );
endmodule
