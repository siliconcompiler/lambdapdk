// //#############################################################################
// //# Function: Tie Low Cell                                                    #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_tielo #(
//     parameter PROP = "DEFAULT"
// ) (
//     output z
// );
// 
//   assign z = 1'b0;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_tielo.v:10.1-18.10" *)
module la_tielo (
    z
);
  (* src = "inputs/la_tielo.v:13.12-13.13" *)
  output z;
  wire z;
  TIELOx1_ASAP7_75t_L _0_ (.L(z));
endmodule
