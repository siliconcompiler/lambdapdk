// //#############################################################################
// //# Function: Or-And-Inverter (oai221) Gate                                   #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_oai221 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a0,
//     input  a1,
//     input  b0,
//     input  b1,
//     input  c0,
//     output z
// );
// 
//   assign z = ~((a0 | a1) & (b0 | b1) & (c0));
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_oai221.v:10.1-23.10" *)
module la_oai221 (
    a0,
    a1,
    b0,
    b1,
    c0,
    z
);
  (* src = "inputs/la_oai221.v:13.12-13.14" *)
  input a0;
  wire a0;
  (* src = "inputs/la_oai221.v:14.12-14.14" *)
  input a1;
  wire a1;
  (* src = "inputs/la_oai221.v:15.12-15.14" *)
  input b0;
  wire b0;
  (* src = "inputs/la_oai221.v:16.12-16.14" *)
  input b1;
  wire b1;
  (* src = "inputs/la_oai221.v:17.12-17.14" *)
  input c0;
  wire c0;
  (* src = "inputs/la_oai221.v:18.12-18.13" *)
  output z;
  wire z;
  sky130_fd_sc_hd__o221ai_4 _0_ (
      .A1(a1),
      .A2(a0),
      .B1(b1),
      .B2(b0),
      .C1(c0),
      .Y (z)
  );
endmodule
