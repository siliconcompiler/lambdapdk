// //#############################################################################
// //# Function: Dual data rate input buffer                                     #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_iddr #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      clk,      // clock
//     input      in,       // data input sampled on both edges of clock
//     output reg outrise,  // rising edge sample
//     output reg outfall   // falling edge sample
// );
// 
//   // Negedge Sample
//   always @(negedge clk) outfall <= in;
// 
//   // Posedge Sample
//   reg inrise;
//   always @(posedge clk) inrise <= in;
// 
//   // Posedge Latch (for hold)
//   always @(clk or inrise) if (~clk) outrise <= inrise;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_iddr.v:10.1-29.10" *)
module la_iddr (
    clk,
    in,
    outrise,
    outfall
);
  wire _0_;
  wire _1_;
  (* src = "inputs/la_iddr.v:13.16-13.19" *)
  input clk;
  wire clk;
  (* src = "inputs/la_iddr.v:14.16-14.18" *)
  input in;
  wire in;
  (* src = "inputs/la_iddr.v:23.7-23.13" *)
  wire inrise;
  (* src = "inputs/la_iddr.v:16.16-16.23" *)
  output outfall;
  wire outfall;
  (* src = "inputs/la_iddr.v:15.16-15.23" *)
  output outrise;
  wire outrise;
  INVx2_ASAP7_75t_SL _2_ (
      .A(_0_),
      .Y(outfall)
  );
  INVx2_ASAP7_75t_SL _3_ (
      .A(_1_),
      .Y(inrise)
  );
  (* module_not_derived = 32'b00000000000000000000000000000001 *)
      (* src = "inputs/la_iddr.v:27.3-27.55|/home/pgadfort/lambdapdk/lambdapdk/asap7/libs/asap7sc7p5t_slvt/techmap/yosys/cells_latch.v:10.24-14.10" *)
  DLLx1_ASAP7_75t_SL _4_ (
      .CLK(clk),
      .D  (inrise),
      .Q  (outrise)
  );
  (* src = "inputs/la_iddr.v:24.3-24.38" *)
  DFFHQNx1_ASAP7_75t_SL _5_ (
      .CLK(clk),
      .D  (in),
      .QN (_1_)
  );
  (* src = "inputs/la_iddr.v:20.3-20.39" *)
  DFFLQNx1_ASAP7_75t_SL _6_ (
      .CLK(clk),
      .D  (in),
      .QN (_0_)
  );
endmodule
