VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

SITE IO_CORNER_75X75
  CLASS PAD ;
  SIZE 75.000 BY 75.000 ;
END IO_CORNER_75X75

SITE IO_SITE_75_H
  CLASS PAD ;
  SIZE 75.000 BY 1.000 ;
END IO_SITE_75_H

SITE IO_SITE_75_V
  CLASS PAD ;
  SIZE 1.000 BY 75.000 ;
END IO_SITE_75_V

MACRO FAKEIO7_BIDIR_V
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 40.000 BY 75.000 ;
  SITE IO_SITE_75_V ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Pad ;
      RECT 10.000 65.000 30.000 70.000 ;
    END
  END PAD
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 55.000 40.000 60.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 45.000 40.000 50.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 35.000 40.000 40.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 25.000 40.000 30.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 19.000 40.000 21.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 15.000 40.000 17.000 ;
    END
  END RING[1]
  PIN IN_ENABLE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
      RECT 4.968 0.000 4.986 1.000 ;
    END
  END IN_ENABLE
  PIN OUT_ENABLE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
      RECT 5.328 0.000 5.346 1.000 ;
    END
  END OUT_ENABLE
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
      RECT 5.688 0.000 5.706 1.000 ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
      RECT 6.048 0.000 6.066 1.000 ;
    END
  END Z
  PIN PULLDOWN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
      RECT 6.408 0.000 6.426 1.000 ;
    END
  END PULLDOWN
  PIN PULLUP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
      RECT 6.768 0.000 6.786 1.000 ;
    END
  END PULLUP
  PIN DRIVE0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
      RECT 6.768 0.000 6.786 1.000 ;
    END
  END DRIVE0
  PIN DRIVE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
      RECT 7.128 0.000 7.146 1.000 ;
    END
  END DRIVE1
  OBS
    LAYER M1 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V1 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M2 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V2 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M3 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V3 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M4 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V4 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M5 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V5 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M6 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V6 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M7 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V7 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M8 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V8 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M9 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V9 ;
    RECT  0.000 0.000 40.000 75.000 ;
  END
END FAKEIO7_BIDIR_V

MACRO FAKEIO7_POC_V
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 10.000 BY 75.000 ;
  SITE IO_SITE_75_V ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 55.000 10.000 60.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 45.000 10.000 50.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 35.000 10.000 40.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 25.000 10.000 30.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 19.000 10.000 21.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 15.000 10.000 17.000 ;
    END
  END RING[1]
  PIN MODE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
      RECT 4.968 0.000 4.986 1.000 ;
    END
  END MODE
  OBS
    LAYER M1 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER V1 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER M2 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER V2 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER M3 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER V3 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER M4 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER V4 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER M5 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER V5 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER M6 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER V6 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER M7 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER V7 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER M8 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER V8 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER M9 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER V9 ;
    RECT  0.000 0.000 10.000 75.000 ;
  END
END FAKEIO7_POC_V

MACRO FAKEIO7_DVDD_V
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 40.000 BY 75.000 ;
  SITE IO_SITE_75_V ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 55.000 40.000 60.000 ;
    END
    PORT
      LAYER Pad ;
      RECT 10.000 65.000 30.000 70.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 45.000 40.000 50.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 35.000 40.000 40.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 25.000 40.000 30.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 19.000 40.000 21.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 15.000 40.000 17.000 ;
    END
  END RING[1]
  OBS
    LAYER M1 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V1 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M2 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V2 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M3 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V3 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M4 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V4 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M5 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V5 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M6 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V6 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M7 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V7 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M8 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V8 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M9 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V9 ;
    RECT  0.000 0.000 40.000 75.000 ;
  END
END FAKEIO7_DVDD_V

MACRO FAKEIO7_DVSS_V
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 40.000 BY 75.000 ;
  SITE IO_SITE_75_V ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 55.000 40.000 60.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 45.000 40.000 50.000 ;
    END
    PORT
      LAYER Pad ;
      RECT 10.000 65.000 30.000 70.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 35.000 40.000 40.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 25.000 40.000 30.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 19.000 40.000 21.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 15.000 40.000 17.000 ;
    END
  END RING[1]
  OBS
    LAYER M1 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V1 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M2 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V2 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M3 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V3 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M4 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V4 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M5 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V5 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M6 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V6 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M7 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V7 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M8 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V8 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M9 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V9 ;
    RECT  0.000 0.000 40.000 75.000 ;
  END
END FAKEIO7_DVSS_V

MACRO FAKEIO7_VDDCLAMP_V
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 40.000 BY 75.000 ;
  SITE IO_SITE_75_V ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 55.000 40.000 60.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 45.000 40.000 50.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 35.000 40.000 40.000 ;
    END
  END VDD
  PIN VDDCLAMP
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Pad ;
      RECT 10.000 65.000 30.000 70.000 ;
    END
    PORT
      LAYER M5 ;
      RECT 10.000 0.000 30.000 2.000 ;
      LAYER M6 ;
      RECT 10.000 0.000 30.000 2.000 ;
      LAYER M7 ;
      RECT 10.000 0.000 30.000 2.000 ;
      LAYER M8 ;
      RECT 10.000 0.000 30.000 2.000 ;
      LAYER M9 ;
      RECT 10.000 0.000 30.000 2.000 ;
    END
  END VDDCLAMP
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 25.000 40.000 30.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 19.000 40.000 21.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 15.000 40.000 17.000 ;
    END
  END RING[1]
  OBS
    LAYER M1 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V1 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M2 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V2 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M3 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V3 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M4 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V4 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M5 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V5 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M6 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V6 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M7 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V7 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M8 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V8 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M9 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V9 ;
    RECT  0.000 0.000 40.000 75.000 ;
  END
END FAKEIO7_VDDCLAMP_V

MACRO FAKEIO7_VDD_V
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 40.000 BY 75.000 ;
  SITE IO_SITE_75_V ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 55.000 40.000 60.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 45.000 40.000 50.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 35.000 40.000 40.000 ;
    END
    PORT
      LAYER Pad ;
      RECT 10.000 65.000 30.000 70.000 ;
    END
    PORT
      LAYER M5 ;
      RECT 10.000 0.000 30.000 2.000 ;
      LAYER M6 ;
      RECT 10.000 0.000 30.000 2.000 ;
      LAYER M7 ;
      RECT 10.000 0.000 30.000 2.000 ;
      LAYER M8 ;
      RECT 10.000 0.000 30.000 2.000 ;
      LAYER M9 ;
      RECT 10.000 0.000 30.000 2.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 25.000 40.000 30.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 19.000 40.000 21.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 15.000 40.000 17.000 ;
    END
  END RING[1]
  OBS
    LAYER M1 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V1 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M2 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V2 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M3 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V3 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M4 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V4 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M5 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V5 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M6 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V6 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M7 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V7 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M8 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V8 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M9 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V9 ;
    RECT  0.000 0.000 40.000 75.000 ;
  END
END FAKEIO7_VDD_V

MACRO FAKEIO7_VSS_V
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 40.000 BY 75.000 ;
  SITE IO_SITE_75_V ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 55.000 40.000 60.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 45.000 40.000 50.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 35.000 40.000 40.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 25.000 40.000 30.000 ;
    END
    PORT
      LAYER Pad ;
      RECT 10.000 65.000 30.000 70.000 ;
    END
    PORT
      LAYER M5 ;
      RECT 10.000 0.000 30.000 2.000 ;
      LAYER M6 ;
      RECT 10.000 0.000 30.000 2.000 ;
      LAYER M7 ;
      RECT 10.000 0.000 30.000 2.000 ;
      LAYER M8 ;
      RECT 10.000 0.000 30.000 2.000 ;
      LAYER M9 ;
      RECT 10.000 0.000 30.000 2.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 19.000 40.000 21.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 15.000 40.000 17.000 ;
    END
  END RING[1]
  OBS
    LAYER M1 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V1 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M2 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V2 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M3 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V3 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M4 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V4 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M5 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V5 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M6 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V6 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M7 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V7 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M8 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V8 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M9 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V9 ;
    RECT  0.000 0.000 40.000 75.000 ;
  END
END FAKEIO7_VSS_V

MACRO FAKEIO7_ANALOG_V
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 40.000 BY 75.000 ;
  SITE IO_SITE_75_V ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Pad ;
      RECT 10.000 65.000 30.000 70.000 ;
    END
  END PAD
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 55.000 40.000 60.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 45.000 40.000 50.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 35.000 40.000 40.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 25.000 40.000 30.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 19.000 40.000 21.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 15.000 40.000 17.000 ;
    END
  END RING[1]
  PIN AIO[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
      RECT 4.968 0.000 4.986 1.000 ;
    END
  END AIO[0]
  PIN AIO[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
      RECT 5.328 0.000 5.346 1.000 ;
    END
  END AIO[1]
  PIN AIO[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
      RECT 5.688 0.000 5.706 1.000 ;
    END
  END AIO[2]
  OBS
    LAYER M1 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V1 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M2 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V2 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M3 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V3 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M4 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V4 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M5 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V5 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M6 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V6 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M7 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V7 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M8 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V8 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER M9 ;
    RECT  0.000 0.000 40.000 75.000 ;
    LAYER V9 ;
    RECT  0.000 0.000 40.000 75.000 ;
  END
END FAKEIO7_ANALOG_V

MACRO FAKEIO7_FILL1_V
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 1.000 BY 75.000 ;
  SITE IO_SITE_75_V ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 55.000 1.000 60.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 45.000 1.000 50.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 35.000 1.000 40.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 25.000 1.000 30.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 19.000 1.000 21.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 15.000 1.000 17.000 ;
    END
  END RING[1]
  OBS
    LAYER M1 ;
    RECT  0.000 0.000 1.000 75.000 ;
    LAYER V1 ;
    RECT  0.000 0.000 1.000 75.000 ;
    LAYER M2 ;
    RECT  0.000 0.000 1.000 75.000 ;
    LAYER V2 ;
    RECT  0.000 0.000 1.000 75.000 ;
    LAYER M3 ;
    RECT  0.000 0.000 1.000 75.000 ;
    LAYER V3 ;
    RECT  0.000 0.000 1.000 75.000 ;
    LAYER M4 ;
    RECT  0.000 0.000 1.000 75.000 ;
    LAYER V4 ;
    RECT  0.000 0.000 1.000 75.000 ;
    LAYER M5 ;
    RECT  0.000 0.000 1.000 75.000 ;
    LAYER V5 ;
    RECT  0.000 0.000 1.000 75.000 ;
    LAYER M6 ;
    RECT  0.000 0.000 1.000 75.000 ;
    LAYER V6 ;
    RECT  0.000 0.000 1.000 75.000 ;
    LAYER M7 ;
    RECT  0.000 0.000 1.000 75.000 ;
    LAYER V7 ;
    RECT  0.000 0.000 1.000 75.000 ;
    LAYER M8 ;
    RECT  0.000 0.000 1.000 75.000 ;
    LAYER V8 ;
    RECT  0.000 0.000 1.000 75.000 ;
    LAYER M9 ;
    RECT  0.000 0.000 1.000 75.000 ;
    LAYER V9 ;
    RECT  0.000 0.000 1.000 75.000 ;
  END
END FAKEIO7_FILL1_V

MACRO FAKEIO7_FILL5_V
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 5.000 BY 75.000 ;
  SITE IO_SITE_75_V ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 55.000 5.000 60.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 45.000 5.000 50.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 35.000 5.000 40.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 25.000 5.000 30.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 19.000 5.000 21.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 15.000 5.000 17.000 ;
    END
  END RING[1]
  OBS
    LAYER M1 ;
    RECT  0.000 0.000 5.000 75.000 ;
    LAYER V1 ;
    RECT  0.000 0.000 5.000 75.000 ;
    LAYER M2 ;
    RECT  0.000 0.000 5.000 75.000 ;
    LAYER V2 ;
    RECT  0.000 0.000 5.000 75.000 ;
    LAYER M3 ;
    RECT  0.000 0.000 5.000 75.000 ;
    LAYER V3 ;
    RECT  0.000 0.000 5.000 75.000 ;
    LAYER M4 ;
    RECT  0.000 0.000 5.000 75.000 ;
    LAYER V4 ;
    RECT  0.000 0.000 5.000 75.000 ;
    LAYER M5 ;
    RECT  0.000 0.000 5.000 75.000 ;
    LAYER V5 ;
    RECT  0.000 0.000 5.000 75.000 ;
    LAYER M6 ;
    RECT  0.000 0.000 5.000 75.000 ;
    LAYER V6 ;
    RECT  0.000 0.000 5.000 75.000 ;
    LAYER M7 ;
    RECT  0.000 0.000 5.000 75.000 ;
    LAYER V7 ;
    RECT  0.000 0.000 5.000 75.000 ;
    LAYER M8 ;
    RECT  0.000 0.000 5.000 75.000 ;
    LAYER V8 ;
    RECT  0.000 0.000 5.000 75.000 ;
    LAYER M9 ;
    RECT  0.000 0.000 5.000 75.000 ;
    LAYER V9 ;
    RECT  0.000 0.000 5.000 75.000 ;
  END
END FAKEIO7_FILL5_V

MACRO FAKEIO7_FILL10_V
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 10.000 BY 75.000 ;
  SITE IO_SITE_75_V ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 55.000 10.000 60.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 45.000 10.000 50.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 35.000 10.000 40.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 25.000 10.000 30.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 19.000 10.000 21.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 15.000 10.000 17.000 ;
    END
  END RING[1]
  OBS
    LAYER M1 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER V1 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER M2 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER V2 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER M3 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER V3 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER M4 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER V4 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER M5 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER V5 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER M6 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER V6 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER M7 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER V7 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER M8 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER V8 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER M9 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER V9 ;
    RECT  0.000 0.000 10.000 75.000 ;
  END
END FAKEIO7_FILL10_V

MACRO FAKEIO7_FILL20_V
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 20.000 BY 75.000 ;
  SITE IO_SITE_75_V ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 55.000 20.000 60.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 45.000 20.000 50.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 35.000 20.000 40.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 25.000 20.000 30.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 19.000 20.000 21.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 15.000 20.000 17.000 ;
    END
  END RING[1]
  OBS
    LAYER M1 ;
    RECT  0.000 0.000 20.000 75.000 ;
    LAYER V1 ;
    RECT  0.000 0.000 20.000 75.000 ;
    LAYER M2 ;
    RECT  0.000 0.000 20.000 75.000 ;
    LAYER V2 ;
    RECT  0.000 0.000 20.000 75.000 ;
    LAYER M3 ;
    RECT  0.000 0.000 20.000 75.000 ;
    LAYER V3 ;
    RECT  0.000 0.000 20.000 75.000 ;
    LAYER M4 ;
    RECT  0.000 0.000 20.000 75.000 ;
    LAYER V4 ;
    RECT  0.000 0.000 20.000 75.000 ;
    LAYER M5 ;
    RECT  0.000 0.000 20.000 75.000 ;
    LAYER V5 ;
    RECT  0.000 0.000 20.000 75.000 ;
    LAYER M6 ;
    RECT  0.000 0.000 20.000 75.000 ;
    LAYER V6 ;
    RECT  0.000 0.000 20.000 75.000 ;
    LAYER M7 ;
    RECT  0.000 0.000 20.000 75.000 ;
    LAYER V7 ;
    RECT  0.000 0.000 20.000 75.000 ;
    LAYER M8 ;
    RECT  0.000 0.000 20.000 75.000 ;
    LAYER V8 ;
    RECT  0.000 0.000 20.000 75.000 ;
    LAYER M9 ;
    RECT  0.000 0.000 20.000 75.000 ;
    LAYER V9 ;
    RECT  0.000 0.000 20.000 75.000 ;
  END
END FAKEIO7_FILL20_V

MACRO FAKEIO7_BREAKER_V
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 10.000 BY 75.000 ;
  SITE IO_SITE_75_V ;
  PIN DVDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 55.000 3.000 60.000 ;
    END
  END DVDDA
  PIN DVDDB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 7.000 55.000 10.000 60.000 ;
    END
  END DVDDB
  PIN DVSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 45.000 3.000 50.000 ;
    END
  END DVSSA
  PIN DVSSB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 7.000 45.000 10.000 50.000 ;
    END
  END DVSSB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 35.000 3.000 40.000 ;
    END
  END VDDA
  PIN VDDB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 7.000 35.000 10.000 40.000 ;
    END
  END VDDB
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 25.000 10.000 30.000 ;
    END
  END VSS
  PIN RINGA[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 19.000 3.000 21.000 ;
    END
  END RINGA[0]
  PIN RINGB[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 7.000 19.000 10.000 21.000 ;
    END
  END RINGB[0]
  PIN RINGA[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 15.000 3.000 17.000 ;
    END
  END RINGA[1]
  PIN RINGB[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 7.000 15.000 10.000 17.000 ;
    END
  END RINGB[1]
  OBS
    LAYER M1 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER V1 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER M2 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER V2 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER M3 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER V3 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER M4 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER V4 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER M5 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER V5 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER M6 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER V6 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER M7 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER V7 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER M8 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER V8 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER M9 ;
    RECT  0.000 0.000 10.000 75.000 ;
    LAYER V9 ;
    RECT  0.000 0.000 10.000 75.000 ;
  END
END FAKEIO7_BREAKER_V

MACRO FAKEIO7_DIFFTX_V
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 80.000 BY 75.000 ;
  SITE IO_SITE_75_V ;
  PIN PADP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Pad ;
      RECT 10.000 65.000 30.000 70.000 ;
    END
  END PADP
  PIN PADN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Pad ;
      RECT 50.000 65.000 70.000 70.000 ;
    END
  END PADN
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 55.000 80.000 60.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 45.000 80.000 50.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 35.000 80.000 40.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 25.000 80.000 30.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 19.000 80.000 21.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 15.000 80.000 17.000 ;
    END
  END RING[1]
  PIN OUT_ENABLE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
      RECT 5.328 0.000 5.346 1.000 ;
    END
  END OUT_ENABLE
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
      RECT 5.688 0.000 5.706 1.000 ;
    END
  END A
  PIN DRIVE0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
      RECT 6.768 0.000 6.786 1.000 ;
    END
  END DRIVE0
  PIN DRIVE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
      RECT 7.128 0.000 7.146 1.000 ;
    END
  END DRIVE1
  OBS
    LAYER M1 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER V1 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER M2 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER V2 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER M3 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER V3 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER M4 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER V4 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER M5 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER V5 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER M6 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER V6 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER M7 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER V7 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER M8 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER V8 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER M9 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER V9 ;
    RECT  0.000 0.000 80.000 75.000 ;
  END
END FAKEIO7_DIFFTX_V

MACRO FAKEIO7_DIFFRX_V
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 80.000 BY 75.000 ;
  SITE IO_SITE_75_V ;
  PIN PADP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Pad ;
      RECT 10.000 65.000 30.000 70.000 ;
    END
  END PADP
  PIN PADN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Pad ;
      RECT 50.000 65.000 70.000 70.000 ;
    END
  END PADN
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 55.000 80.000 60.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 45.000 80.000 50.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 35.000 80.000 40.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 25.000 80.000 30.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 19.000 80.000 21.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 15.000 80.000 17.000 ;
    END
  END RING[1]
  PIN IN_ENABLE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
      RECT 4.968 0.000 4.986 1.000 ;
    END
  END IN_ENABLE
  PIN ZP
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
      RECT 5.688 0.000 5.706 1.000 ;
    END
  END ZP
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
      RECT 6.048 0.000 6.066 1.000 ;
    END
  END ZN
  PIN PULLDOWN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
      RECT 6.408 0.000 6.426 1.000 ;
    END
  END PULLDOWN
  PIN PULLUP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
      RECT 6.768 0.000 6.786 1.000 ;
    END
  END PULLUP
  OBS
    LAYER M1 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER V1 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER M2 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER V2 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER M3 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER V3 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER M4 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER V4 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER M5 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER V5 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER M6 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER V6 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER M7 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER V7 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER M8 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER V8 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER M9 ;
    RECT  0.000 0.000 80.000 75.000 ;
    LAYER V9 ;
    RECT  0.000 0.000 80.000 75.000 ;
  END
END FAKEIO7_DIFFRX_V

MACRO FAKEIO7_CORNER
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 75.000 BY 75.000 ;
  SITE IO_CORNER_75X75 ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 55.000 3.000 60.000 ;
    END
    PORT
      LAYER M9 ;
      RECT 55.000 0.000 60.000 3.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 45.000 3.000 50.000 ;
    END
    PORT
      LAYER M9 ;
      RECT 45.000 0.000 50.000 3.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 0.000 35.000 3.000 40.000 ;
    END
    PORT
      LAYER M9 ;
      RECT 35.000 0.000 40.000 3.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 0.000 25.000 3.000 30.000 ;
    END
    PORT
      LAYER M9 ;
      RECT 25.000 0.000 30.000 3.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 19.000 3.000 21.000 ;
    END
    PORT
      LAYER M8 ;
      RECT 19.000 0.000 21.000 3.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 0.000 15.000 3.000 17.000 ;
    END
    PORT
      LAYER M8 ;
      RECT 15.000 0.000 17.000 3.000 ;
    END
  END RING[1]
  OBS
    LAYER M1 ;
    RECT  0.000 0.000 75.000 75.000 ;
    LAYER V1 ;
    RECT  0.000 0.000 75.000 75.000 ;
    LAYER M2 ;
    RECT  0.000 0.000 75.000 75.000 ;
    LAYER V2 ;
    RECT  0.000 0.000 75.000 75.000 ;
    LAYER M3 ;
    RECT  0.000 0.000 75.000 75.000 ;
    LAYER V3 ;
    RECT  0.000 0.000 75.000 75.000 ;
    LAYER M4 ;
    RECT  0.000 0.000 75.000 75.000 ;
    LAYER V4 ;
    RECT  0.000 0.000 75.000 75.000 ;
    LAYER M5 ;
    RECT  0.000 0.000 75.000 75.000 ;
    LAYER V5 ;
    RECT  0.000 0.000 75.000 75.000 ;
    LAYER M6 ;
    RECT  0.000 0.000 75.000 75.000 ;
    LAYER V6 ;
    RECT  0.000 0.000 75.000 75.000 ;
    LAYER M7 ;
    RECT  0.000 0.000 75.000 75.000 ;
    LAYER V7 ;
    RECT  0.000 0.000 75.000 75.000 ;
    LAYER M8 ;
    RECT  0.000 0.000 75.000 75.000 ;
    LAYER V8 ;
    RECT  0.000 0.000 75.000 75.000 ;
    LAYER M9 ;
    RECT  0.000 0.000 75.000 75.000 ;
    LAYER V9 ;
    RECT  0.000 0.000 75.000 75.000 ;
  END
END FAKEIO7_CORNER

MACRO FAKEIO7_BUMP_SMALL
  CLASS COVER BUMP ;
  SYMMETRY X Y R90 ;
  SIZE 30.000 BY 30.000 ;
  ORIGIN 15.000 15.000 ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Pad ;
      POLYGON -6.213 -15.000 -15.000 -6.213 -15.000 6.213 -6.213 15.000 6.213 15.000 15.000 6.213 15.000 -6.213 6.213 -15.000 ;
    END
  END PAD
  OBS
    LAYER V9 ;
    POLYGON -6.213 -15.000 -15.000 -6.213 -15.000 6.213 -6.213 15.000 6.213 15.000 15.000 6.213 15.000 -6.213 6.213 -15.000 ;
  END
END FAKEIO7_BUMP_SMALL

MACRO FAKEIO7_BUMP_LARGE
  CLASS COVER BUMP ;
  SYMMETRY X Y R90 ;
  SIZE 50.000 BY 50.000 ;
  ORIGIN 25.000 25.000 ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Pad ;
      POLYGON -10.355 -25.000 -25.000 -10.355 -25.000 10.355 -10.355 25.000 10.355 25.000 25.000 10.355 25.000 -10.355 10.355 -25.000 ;
    END
  END PAD
  OBS
    LAYER V9 ;
    POLYGON -9.113 -22.000  -22.000 -9.113  -22.000 9.113 -9.113 22.000 9.113 22.000 22.000 9.113 22.000 -9.113 9.113 -22.000 ;
  END
END FAKEIO7_BUMP_LARGE

MACRO FAKEIO7_BIDIR_H
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 75.000 BY 40.000 ;
  SITE IO_SITE_75_H ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Pad ;
      RECT 65.000 10.000 70.000 30.000 ;
    END
  END PAD
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 55.000 0.000 60.000 40.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 45.000 0.000 50.000 40.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 35.000 0.000 40.000 40.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 25.000 0.000 30.000 40.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 19.000 0.000 21.000 40.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 15.000 0.000 17.000 40.000 ;
    END
  END RING[1]
  PIN IN_ENABLE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.968 1.000 4.986 ;
    END
  END IN_ENABLE
  PIN OUT_ENABLE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.328 1.000 5.346 ;
    END
  END OUT_ENABLE
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.688 1.000 5.706 ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.048 1.000 6.066 ;
    END
  END Z
  PIN PULLDOWN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.408 1.000 6.426 ;
    END
  END PULLDOWN
  PIN PULLUP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.768 1.000 6.786 ;
    END
  END PULLUP
  PIN DRIVE0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.768 1.000 6.786 ;
    END
  END DRIVE0
  PIN DRIVE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.128 1.000 7.146 ;
    END
  END DRIVE1
  OBS
    LAYER M1 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V1 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M2 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V2 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M3 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V3 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M4 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V4 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M5 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V5 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M6 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V6 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M7 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V7 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M8 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V8 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M9 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V9 ;
    RECT 0.000 0.000 75.000 40.000 ;
  END
END FAKEIO7_BIDIR_H

MACRO FAKEIO7_POC_H
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 75.000 BY 10.000 ;
  SITE IO_SITE_75_H ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 55.000 0.000 60.000 10.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 45.000 0.000 50.000 10.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 35.000 0.000 40.000 10.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 25.000 0.000 30.000 10.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 19.000 0.000 21.000 10.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 15.000 0.000 17.000 10.000 ;
    END
  END RING[1]
  PIN MODE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.968 1.000 4.986 ;
    END
  END MODE
  OBS
    LAYER M1 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER V1 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER M2 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER V2 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER M3 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER V3 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER M4 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER V4 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER M5 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER V5 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER M6 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER V6 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER M7 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER V7 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER M8 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER V8 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER M9 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER V9 ;
    RECT 0.000 0.000 75.000 10.000 ;
  END
END FAKEIO7_POC_H

MACRO FAKEIO7_DVDD_H
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 75.000 BY 40.000 ;
  SITE IO_SITE_75_H ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 55.000 0.000 60.000 40.000 ;
    END
    PORT
      LAYER Pad ;
      RECT 65.000 10.000 70.000 30.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 45.000 0.000 50.000 40.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 35.000 0.000 40.000 40.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 25.000 0.000 30.000 40.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 19.000 0.000 21.000 40.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 15.000 0.000 17.000 40.000 ;
    END
  END RING[1]
  OBS
    LAYER M1 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V1 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M2 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V2 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M3 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V3 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M4 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V4 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M5 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V5 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M6 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V6 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M7 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V7 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M8 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V8 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M9 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V9 ;
    RECT 0.000 0.000 75.000 40.000 ;
  END
END FAKEIO7_DVDD_H

MACRO FAKEIO7_DVSS_H
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 75.000 BY 40.000 ;
  SITE IO_SITE_75_H ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 55.000 0.000 60.000 40.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 45.000 0.000 50.000 40.000 ;
    END
    PORT
      LAYER Pad ;
      RECT 65.000 10.000 70.000 30.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 35.000 0.000 40.000 40.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 25.000 0.000 30.000 40.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 19.000 0.000 21.000 40.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 15.000 0.000 17.000 40.000 ;
    END
  END RING[1]
  OBS
    LAYER M1 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V1 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M2 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V2 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M3 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V3 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M4 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V4 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M5 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V5 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M6 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V6 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M7 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V7 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M8 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V8 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M9 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V9 ;
    RECT 0.000 0.000 75.000 40.000 ;
  END
END FAKEIO7_DVSS_H

MACRO FAKEIO7_VDD_H
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 75.000 BY 40.000 ;
  SITE IO_SITE_75_H ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 55.000 0.000 60.000 40.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 45.000 0.000 50.000 40.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 35.000 0.000 40.000 40.000 ;
    END
    PORT
      LAYER Pad ;
      RECT 65.000 10.000 70.000 30.000 ;
    END
    PORT
      LAYER M5 ;
      RECT 0.000 10.000 2.000 30.000 ;
      LAYER M6 ;
      RECT 0.000 10.000 2.000 30.000 ;
      LAYER M7 ;
      RECT 0.000 10.000 2.000 30.000 ;
      LAYER M8 ;
      RECT 0.000 10.000 2.000 30.000 ;
      LAYER M9 ;
      RECT 0.000 10.000 2.000 30.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 25.000 0.000 30.000 40.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 19.000 0.000 21.000 40.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 15.000 0.000 17.000 40.000 ;
    END
  END RING[1]
  OBS
    LAYER M1 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V1 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M2 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V2 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M3 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V3 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M4 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V4 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M5 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V5 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M6 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V6 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M7 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V7 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M8 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V8 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M9 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V9 ;
    RECT 0.000 0.000 75.000 40.000 ;
  END
END FAKEIO7_VDD_H

MACRO FAKEIO7_VSS_H
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 75.000 BY 40.000 ;
  SITE IO_SITE_75_H ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 55.000 0.000 60.000 40.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 45.000 0.000 50.000 40.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 35.000 0.000 40.000 40.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 25.000 0.000 30.000 40.000 ;
    END
    PORT
      LAYER Pad ;
      RECT 65.000 10.000 70.000 30.000 ;
    END
    PORT
      LAYER M5 ;
      RECT 0.000 10.000 2.000 30.000 ;
      LAYER M6 ;
      RECT 0.000 10.000 2.000 30.000 ;
      LAYER M7 ;
      RECT 0.000 10.000 2.000 30.000 ;
      LAYER M8 ;
      RECT 0.000 10.000 2.000 30.000 ;
      LAYER M9 ;
      RECT 0.000 10.000 2.000 30.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 19.000 0.000 21.000 40.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 15.000 0.000 17.000 40.000 ;
    END
  END RING[1]
  OBS
    LAYER M1 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V1 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M2 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V2 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M3 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V3 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M4 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V4 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M5 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V5 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M6 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V6 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M7 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V7 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M8 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V8 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M9 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V9 ;
    RECT 0.000 0.000 75.000 40.000 ;
  END
END FAKEIO7_VSS_H

MACRO FAKEIO7_ANALOG_H
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 75.000 BY 40.000 ;
  SITE IO_SITE_75_H ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Pad ;
      RECT 65.000 10.000 70.000 30.000 ;
    END
  END PAD
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 55.000 0.000 60.000 40.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 45.000 0.000 50.000 40.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 35.000 0.000 40.000 40.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 25.000 0.000 30.000 40.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 19.000 0.000 21.000 40.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 15.000 0.000 17.000 40.000 ;
    END
  END RING[1]
  PIN AIO[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.968 1.000 4.986 ;
    END
  END AIO[0]
  PIN AIO[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.328 1.000 5.346 ;
    END
  END AIO[1]
  PIN AIO[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.688 1.000 5.706 ;
    END
  END AIO[2]
  OBS
    LAYER M1 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V1 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M2 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V2 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M3 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V3 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M4 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V4 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M5 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V5 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M6 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V6 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M7 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V7 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M8 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V8 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M9 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V9 ;
    RECT 0.000 0.000 75.000 40.000 ;
  END
END FAKEIO7_ANALOG_H

MACRO FAKEIO7_FILL1_H
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 75.000 BY 1.000 ;
  SITE IO_SITE_75_H ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 55.000 0.000 60.000 1.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 45.000 0.000 50.000 1.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 35.000 0.000 40.000 1.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 25.000 0.000 30.000 1.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 19.000 0.000 21.000 1.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 15.000 0.000 17.000 1.000 ;
    END
  END RING[1]
  OBS
    LAYER M1 ;
    RECT 0.000 0.000 75.000 1.000 ;
    LAYER V1 ;
    RECT 0.000 0.000 75.000 1.000 ;
    LAYER M2 ;
    RECT 0.000 0.000 75.000 1.000 ;
    LAYER V2 ;
    RECT 0.000 0.000 75.000 1.000 ;
    LAYER M3 ;
    RECT 0.000 0.000 75.000 1.000 ;
    LAYER V3 ;
    RECT 0.000 0.000 75.000 1.000 ;
    LAYER M4 ;
    RECT 0.000 0.000 75.000 1.000 ;
    LAYER V4 ;
    RECT 0.000 0.000 75.000 1.000 ;
    LAYER M5 ;
    RECT 0.000 0.000 75.000 1.000 ;
    LAYER V5 ;
    RECT 0.000 0.000 75.000 1.000 ;
    LAYER M6 ;
    RECT 0.000 0.000 75.000 1.000 ;
    LAYER V6 ;
    RECT 0.000 0.000 75.000 1.000 ;
    LAYER M7 ;
    RECT 0.000 0.000 75.000 1.000 ;
    LAYER V7 ;
    RECT 0.000 0.000 75.000 1.000 ;
    LAYER M8 ;
    RECT 0.000 0.000 75.000 1.000 ;
    LAYER V8 ;
    RECT 0.000 0.000 75.000 1.000 ;
    LAYER M9 ;
    RECT 0.000 0.000 75.000 1.000 ;
    LAYER V9 ;
    RECT 0.000 0.000 75.000 1.000 ;
  END
END FAKEIO7_FILL1_H

MACRO FAKEIO7_FILL5_H
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 75.000 BY 5.000 ;
  SITE IO_SITE_75_H ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 55.000 0.000 60.000 5.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 45.000 0.000 50.000 5.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 35.000 0.000 40.000 5.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 25.000 0.000 30.000 5.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 19.000 0.000 21.000 5.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 15.000 0.000 17.000 5.000 ;
    END
  END RING[1]
  OBS
    LAYER M1 ;
    RECT 0.000 0.000 75.000 5.000 ;
    LAYER V1 ;
    RECT 0.000 0.000 75.000 5.000 ;
    LAYER M2 ;
    RECT 0.000 0.000 75.000 5.000 ;
    LAYER V2 ;
    RECT 0.000 0.000 75.000 5.000 ;
    LAYER M3 ;
    RECT 0.000 0.000 75.000 5.000 ;
    LAYER V3 ;
    RECT 0.000 0.000 75.000 5.000 ;
    LAYER M4 ;
    RECT 0.000 0.000 75.000 5.000 ;
    LAYER V4 ;
    RECT 0.000 0.000 75.000 5.000 ;
    LAYER M5 ;
    RECT 0.000 0.000 75.000 5.000 ;
    LAYER V5 ;
    RECT 0.000 0.000 75.000 5.000 ;
    LAYER M6 ;
    RECT 0.000 0.000 75.000 5.000 ;
    LAYER V6 ;
    RECT 0.000 0.000 75.000 5.000 ;
    LAYER M7 ;
    RECT 0.000 0.000 75.000 5.000 ;
    LAYER V7 ;
    RECT 0.000 0.000 75.000 5.000 ;
    LAYER M8 ;
    RECT 0.000 0.000 75.000 5.000 ;
    LAYER V8 ;
    RECT 0.000 0.000 75.000 5.000 ;
    LAYER M9 ;
    RECT 0.000 0.000 75.000 5.000 ;
    LAYER V9 ;
    RECT 0.000 0.000 75.000 5.000 ;
  END
END FAKEIO7_FILL5_H

MACRO FAKEIO7_FILL10_H
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 75.000 BY 10.000 ;
  SITE IO_SITE_75_H ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 55.000 0.000 60.000 10.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 45.000 0.000 50.000 10.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 35.000 0.000 40.000 10.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 25.000 0.000 30.000 10.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 19.000 0.000 21.000 10.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 15.000 0.000 17.000 10.000 ;
    END
  END RING[1]
  OBS
    LAYER M1 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER V1 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER M2 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER V2 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER M3 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER V3 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER M4 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER V4 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER M5 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER V5 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER M6 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER V6 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER M7 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER V7 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER M8 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER V8 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER M9 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER V9 ;
    RECT 0.000 0.000 75.000 10.000 ;
  END
END FAKEIO7_FILL10_H

MACRO FAKEIO7_FILL20_H
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 75.000 BY 20.000 ;
  SITE IO_SITE_75_H ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 55.000 0.000 60.000 20.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 45.000 0.000 50.000 20.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 35.000 0.000 40.000 20.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 25.000 0.000 30.000 20.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 19.000 0.000 21.000 20.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 15.000 0.000 17.000 20.000 ;
    END
  END RING[1]
  OBS
    LAYER M1 ;
    RECT 0.000 0.000 75.000 20.000 ;
    LAYER V1 ;
    RECT 0.000 0.000 75.000 20.000 ;
    LAYER M2 ;
    RECT 0.000 0.000 75.000 20.000 ;
    LAYER V2 ;
    RECT 0.000 0.000 75.000 20.000 ;
    LAYER M3 ;
    RECT 0.000 0.000 75.000 20.000 ;
    LAYER V3 ;
    RECT 0.000 0.000 75.000 20.000 ;
    LAYER M4 ;
    RECT 0.000 0.000 75.000 20.000 ;
    LAYER V4 ;
    RECT 0.000 0.000 75.000 20.000 ;
    LAYER M5 ;
    RECT 0.000 0.000 75.000 20.000 ;
    LAYER V5 ;
    RECT 0.000 0.000 75.000 20.000 ;
    LAYER M6 ;
    RECT 0.000 0.000 75.000 20.000 ;
    LAYER V6 ;
    RECT 0.000 0.000 75.000 20.000 ;
    LAYER M7 ;
    RECT 0.000 0.000 75.000 20.000 ;
    LAYER V7 ;
    RECT 0.000 0.000 75.000 20.000 ;
    LAYER M8 ;
    RECT 0.000 0.000 75.000 20.000 ;
    LAYER V8 ;
    RECT 0.000 0.000 75.000 20.000 ;
    LAYER M9 ;
    RECT 0.000 0.000 75.000 20.000 ;
    LAYER V9 ;
    RECT 0.000 0.000 75.000 20.000 ;
  END
END FAKEIO7_FILL20_H

MACRO FAKEIO7_BREAKER_H
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 75.000 BY 10.000 ;
  SITE IO_SITE_75_H ;
  PIN DVDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 55.000 0.000 60.000 3.000 ;
    END
  END DVDDA
  PIN DVDDB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 55.000 7.000 60.000 10.000 ;
    END
  END DVDDB
  PIN DVSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 45.000 0.000 50.000 3.000 ;
    END
  END DVSSA
  PIN DVSSB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 45.000 7.000 50.000 10.000 ;
    END
  END DVSSB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 35.000 0.000 40.000 3.000 ;
    END
  END VDDA
  PIN VDDB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 35.000 7.000 40.000 10.000 ;
    END
  END VDDB
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 25.000 0.000 30.000 10.000 ;
    END
  END VSS
  PIN RINGA[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 19.000 0.000 21.000 3.000 ;
    END
  END RINGA[0]
  PIN RINGB[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 19.000 7.000 21.000 10.000 ;
    END
  END RINGB[0]
  PIN RINGA[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 15.000 0.000 17.000 3.000 ;
    END
  END RINGA[1]
  PIN RINGB[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 15.000 7.000 17.000 10.000 ;
    END
  END RINGB[1]
  OBS
    LAYER M1 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER V1 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER M2 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER V2 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER M3 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER V3 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER M4 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER V4 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER M5 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER V5 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER M6 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER V6 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER M7 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER V7 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER M8 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER V8 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER M9 ;
    RECT 0.000 0.000 75.000 10.000 ;
    LAYER V9 ;
    RECT 0.000 0.000 75.000 10.000 ;
  END
END FAKEIO7_BREAKER_H

MACRO FAKEIO7_DIFFTX_H
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 75.000 BY 80.000 ;
  SITE IO_SITE_75_H ;
  PIN PADP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Pad ;
      RECT 65.000 10.000 70.000 30.000 ;
    END
  END PADP
  PIN PADN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Pad ;
      RECT 65.000 50.000 70.000 70.000 ;
    END
  END PADN
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 55.000 0.000 60.000 80.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 45.000 0.000 50.000 80.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 35.000 0.000 40.000 80.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 25.000 0.000 30.000 80.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 19.000 0.000 21.000 80.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 15.000 0.000 17.000 80.000 ;
    END
  END RING[1]
  PIN OUT_ENABLE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.328 1.000 5.346 ;
    END
  END OUT_ENABLE
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.688 1.000 5.706 ;
    END
  END A
  PIN DRIVE0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.768 1.000 6.786 ;
    END
  END DRIVE0
  PIN DRIVE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.128 1.000 7.146 ;
    END
  END DRIVE1
  OBS
    LAYER M1 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER V1 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER M2 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER V2 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER M3 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER V3 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER M4 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER V4 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER M5 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER V5 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER M6 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER V6 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER M7 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER V7 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER M8 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER V8 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER M9 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER V9 ;
    RECT 0.000 0.000 75.000 80.000 ;
  END
END FAKEIO7_DIFFTX_H

MACRO FAKEIO7_DIFFRX_H
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 75.000 BY 80.000 ;
  SITE IO_SITE_75_H ;
  PIN PADP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Pad ;
      RECT 65.000 10.000 70.000 30.000 ;
    END
  END PADP
  PIN PADN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Pad ;
      RECT 65.000 50.000 70.000 70.000 ;
    END
  END PADN
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 55.000 0.000 60.000 80.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 45.000 0.000 50.000 80.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 35.000 0.000 40.000 80.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 25.000 0.000 30.000 80.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 19.000 0.000 21.000 80.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 15.000 0.000 17.000 80.000 ;
    END
  END RING[1]
  PIN IN_ENABLE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.968 1.000 4.986 ;
    END
  END IN_ENABLE
  PIN ZP
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.688 1.000 5.706 ;
    END
  END ZP
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.048 1.000 6.066 ;
    END
  END ZN
  PIN PULLDOWN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.408 1.000 6.426 ;
    END
  END PULLDOWN
  PIN PULLUP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.768 1.000 6.786 ;
    END
  END PULLUP
  OBS
    LAYER M1 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER V1 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER M2 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER V2 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER M3 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER V3 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER M4 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER V4 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER M5 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER V5 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER M6 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER V6 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER M7 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER V7 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER M8 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER V8 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER M9 ;
    RECT 0.000 0.000 75.000 80.000 ;
    LAYER V9 ;
    RECT 0.000 0.000 75.000 80.000 ;
  END
END FAKEIO7_DIFFRX_H

MACRO FAKEIO7_VDDCLAMP_H
  CLASS PAD AREAIO ;
  SYMMETRY X Y ;
  SIZE 75.000 BY 40.000 ;
  SITE IO_SITE_75_H ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 55.000 0.000 60.000 40.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 45.000 0.000 50.000 40.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
      RECT 35.000 0.000 40.000 40.000 ;
    END
  END VDD
  PIN VDDCLAMP
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Pad ;
      RECT 65.000 10.000 70.000 30.000 ;
    END
    PORT
      LAYER M5 ;
      RECT 0.000 10.000 2.000 30.000 ;
      LAYER M6 ;
      RECT 0.000 10.000 2.000 30.000 ;
      LAYER M7 ;
      RECT 0.000 10.000 2.000 30.000 ;
      LAYER M8 ;
      RECT 0.000 10.000 2.000 30.000 ;
      LAYER M9 ;
      RECT 0.000 10.000 2.000 30.000 ;
    END
  END VDDCLAMP
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
      RECT 25.000 0.000 30.000 40.000 ;
    END
  END VSS
  PIN RING[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 19.000 0.000 21.000 40.000 ;
    END
  END RING[0]
  PIN RING[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
      RECT 15.000 0.000 17.000 40.000 ;
    END
  END RING[1]
  OBS
    LAYER M1 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V1 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M2 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V2 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M3 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V3 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M4 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V4 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M5 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V5 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M6 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V6 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M7 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V7 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M8 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V8 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER M9 ;
    RECT 0.000 0.000 75.000 40.000 ;
    LAYER V9 ;
    RECT 0.000 0.000 75.000 40.000 ;
  END
END FAKEIO7_VDDCLAMP_H
