// //#############################################################################
// //# Function:  Positive edge-triggered static D-type flop-flop with async     #
// //#            active low preset.                                             #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_dffsq #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      clk,
//     input      nset,
//     output reg q
// );
// 
//     always @(posedge clk or negedge nset)
//         if (!nset) q <= 1'b1;
//         else q <= d;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
(* keep_hierarchy *)
module la_dffsq (
    d,
    clk,
    nset,
    q
);
  (* src = "generated" *)
  input clk;
  wire clk;
  (* src = "generated" *)
  input d;
  wire d;
  (* src = "generated" *)
  input nset;
  wire nset;
  (* src = "generated" *)
  output q;
  wire q;
  (* src = "generated" *)
  gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 _0_ (
      .CLK(clk),
      .D(d),
      .Q(q),
      .SETN(nset)
  );
endmodule
