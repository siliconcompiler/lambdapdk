// //#############################################################################
// //# Function: And-Or (ao33) Gate                                              #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_ao33 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a0,
//     input  a1,
//     input  a2,
//     input  b0,
//     input  b1,
//     input  b2,
//     output z
// );
// 
//     assign z = (a0 & a1 & a2) | (b0 & b1 & b2);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
(* keep_hierarchy *)
module la_ao33 (
    a0,
    a1,
    a2,
    b0,
    b1,
    b2,
    z
);
  wire _0_;
  wire _1_;
  (* src = "generated" *)
  input a0;
  wire a0;
  (* src = "generated" *)
  input a1;
  wire a1;
  (* src = "generated" *)
  input a2;
  wire a2;
  (* src = "generated" *)
  input b0;
  wire b0;
  (* src = "generated" *)
  input b1;
  wire b1;
  (* src = "generated" *)
  input b2;
  wire b2;
  (* src = "generated" *)
  output z;
  wire z;
  NAND3_X2 _2_ (
      .A1(b2),
      .A2(b1),
      .A3(b0),
      .ZN(_0_)
  );
  NAND3_X2 _3_ (
      .A1(a1),
      .A2(a0),
      .A3(a2),
      .ZN(_1_)
  );
  NAND2_X2 _4_ (
      .A1(_0_),
      .A2(_1_),
      .ZN(z)
  );
endmodule
