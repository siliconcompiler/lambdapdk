// //#############################################################################
// //# Function:  Positive edge-triggered static D-type flop-flop with async     #
// //#            active low reset and scan input                                #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_sdffrq #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      si,
//     input      se,
//     input      clk,
//     input      nreset,
//     output reg q
// );
// 
//     always @(posedge clk or negedge nreset)
//         if (!nreset) q <= 1'b0;
//         else q <= se ? si : d;
// 
// endmodule

/* Generated by Yosys 0.40 (git sha1 a1bb0255d, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_sdffrq(d, si, se, clk, nreset, q);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  input clk;
  wire clk;
  input d;
  wire d;
  input nreset;
  wire nreset;
  output q;
  wire q;
  input se;
  wire se;
  input si;
  wire si;
  INVx1_ASAP7_75t_SL _05_ (
    .A(se),
    .Y(_02_)
  );
  AND2x4_ASAP7_75t_SL _06_ (
    .A(si),
    .B(se),
    .Y(_03_)
  );
  AO21x1_ASAP7_75t_SL _07_ (
    .A1(d),
    .A2(_02_),
    .B(_03_),
    .Y(_00_)
  );
  INVx1_ASAP7_75t_SL _08_ (
    .A(_01_),
    .Y(q)
  );
  DFFASRHQNx1_ASAP7_75t_SL _09_ (
    .CLK(clk),
    .D(_00_),
    .QN(_01_),
    .RESETN(_04_),
    .SETN(nreset)
  );
  TIEHIx1_ASAP7_75t_SL _10_ (
    .H(_04_)
  );
endmodule
