// //#############################################################################
// //# Function: Power isolation circuit                                         #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_isolo #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  iso,  // isolation signal
//     input  in,   // input
//     output out   // out = ~iso & in
// );
// 
//   assign out = ~iso & in;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_isolo.v:10.1-20.10" *)
module la_isolo (
    iso,
    in,
    out
);
  (* src = "inputs/la_isolo.v:14.12-14.14" *)
  input in;
  wire in;
  (* src = "inputs/la_isolo.v:13.12-13.15" *)
  input iso;
  wire iso;
  (* src = "inputs/la_isolo.v:15.12-15.15" *)
  output out;
  wire out;
  sky130_fd_sc_hd__nor2b_4 _0_ (
      .A  (iso),
      .B_N(in),
      .Y  (out)
  );
endmodule
