// Width of padring configuration bus with values
// such as drive strength.

`define LA_PADRING_CFGW n

// Width of ring bus with power, ground, vref signals usually
// connected by abutment in the padring.

`define LA_PADRING_RINGW 8
