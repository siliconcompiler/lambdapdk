// //#############################################################################
// //# Function: Carry Save Adder (3:2)                                          #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_csa32 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     input  b,
//     input  c,
//     output sum,
//     output carry
// );
// 
//     assign sum   = a ^ b ^ c;
//     assign carry = (a & b) | (b & c) | (c & a);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
module la_csa32 (
    a,
    b,
    c,
    sum,
    carry
);
  (* src = "generated" *)
  wire _0_;
  (* src = "generated" *)
  wire _1_;
  (* src = "generated" *)
  input a;
  wire a;
  (* src = "generated" *)
  input b;
  wire b;
  (* src = "generated" *)
  input c;
  wire c;
  (* src = "generated" *)
  output carry;
  wire carry;
  (* src = "generated" *)
  output sum;
  wire sum;
  INVx2_ASAP7_75t_R _2_ (
      .A(_0_),
      .Y(carry)
  );
  INVx2_ASAP7_75t_R _3_ (
      .A(_1_),
      .Y(sum)
  );
  (* module_not_derived = 32'b00000000000000000000000000000001 *) (* src = "generated" *)
  FAx1_ASAP7_75t_R _4_ (
      .A  (a),
      .B  (b),
      .CI (c),
      .CON(_0_),
      .SN (_1_)
  );
endmodule
