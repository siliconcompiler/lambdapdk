// //#############################################################################
// //# Function: 2-Input Clock OR Gate                                           #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_clkor2 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     input  b,
//     output z
// );
// 
//     assign z = a | b;
// 
// endmodule

/* Generated by Yosys 0.40+33 (git sha1 cd1fb8b15, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_clkor2(a, b, z);
  input a;
  wire a;
  input b;
  wire b;
  output z;
  wire z;
  sg13g2_or2_1 _0_ (
    .A(b),
    .B(a),
    .X(z)
  );
endmodule
