// //#############################################################################
// //# Function: Carry Save Adder (4:2) (aka 5:3)                                #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_csa42 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     input  b,
//     input  c,
//     input  d,
//     input  cin,
//     output sum,
//     output carry,
//     output cout
// );
// 
//     assign cout   = (a & b) | (b & c) | (a & c);
//     assign sumint = a ^ b ^ c;
//     assign sum    = cin ^ d ^ sumint;
//     assign carry  = (cin & d) | (cin & sumint) | (d & sumint);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
(* keep_hierarchy *)
module la_csa42 (
    a,
    b,
    c,
    d,
    cin,
    sum,
    carry,
    cout
);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  (* src = "generated" *)
  input a;
  wire a;
  (* src = "generated" *)
  input b;
  wire b;
  (* src = "generated" *)
  input c;
  wire c;
  (* src = "generated" *)
  output carry;
  wire carry;
  (* src = "generated" *)
  input cin;
  wire cin;
  (* src = "generated" *)
  output cout;
  wire cout;
  (* src = "generated" *)
  input d;
  wire d;
  (* src = "generated" *)
  output sum;
  wire sum;
  sky130_fd_sc_hdll__nor2_1 _06_ (
      .A(b),
      .B(a),
      .Y(_05_)
  );
  sky130_fd_sc_hdll__a21oi_1 _07_ (
      .A1(b),
      .A2(a),
      .B1(c),
      .Y (_00_)
  );
  sky130_fd_sc_hdll__nor2_1 _08_ (
      .A(_05_),
      .B(_00_),
      .Y(cout)
  );
  sky130_fd_sc_hdll__xor2_1 _09_ (
      .A(d),
      .B(cin),
      .X(_01_)
  );
  sky130_fd_sc_hdll__xnor3_1 _10_ (
      .A(b),
      .B(a),
      .C(c),
      .X(_02_)
  );
  sky130_fd_sc_hdll__xnor2_2 _11_ (
      .A(_01_),
      .B(_02_),
      .Y(sum)
  );
  sky130_fd_sc_hdll__nand2_6 _12_ (
      .A(d),
      .B(cin),
      .Y(_03_)
  );
  sky130_fd_sc_hdll__nor2_1 _13_ (
      .A(d),
      .B(cin),
      .Y(_04_)
  );
  sky130_fd_sc_hdll__a21oi_2 _14_ (
      .A1(_03_),
      .A2(_02_),
      .B1(_04_),
      .Y (carry)
  );
endmodule
