# Copyright 2024 ZeroASIC Corp
# 
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
# 
#      https://www.apache.org/licenses/LICENSE-2.0
# 
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER metal1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.8 ;
  SPACING 0.4 ;
  WIDTH 0.4 ;
  MAXWIDTH 5.0 ;
END metal1

LAYER via1
  TYPE CUT ;
  SPACING 0.2 ;
  WIDTH 0.2 ;
END via1

LAYER metal2
  TYPE ROUTING ;
  DIRECTION VERITCAL ;
  PITCH 0.8 ;
  SPACING 0.4 ;
  WIDTH 0.4 ;
  MAXWIDTH 5.0 ;
END metal2

LAYER via2
  TYPE CUT ;
  SPACING 0.2 ;
  WIDTH 0.2 ;
END via2

LAYER metal3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.8 ;
  SPACING 0.4 ;
  WIDTH 0.4 ;
  MAXWIDTH 5.0 ;
END metal3

LAYER via3
  TYPE CUT ;
  SPACING 0.2 ;
  WIDTH 0.2 ;
END via3

LAYER topmetal
  TYPE ROUTING ;
  DIRECTION VERITCAL ;
  PITCH 0.8 ;
  SPACING 0.4 ;
  WIDTH 0.4 ;
  MAXWIDTH 5.0 ;
END topmetal

VIA VIA1_1 DEFAULT
  LAYER via1 ;
    RECT -0.100 -0.100 0.100 0.100 ;
  LAYER metal1 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  LAYER metal2 ;
    RECT -0.300 -0.300 0.300 0.300 ;
END VIA1_1

VIA VIA2_1 DEFAULT
  LAYER via2 ;
    RECT -0.100 -0.100 0.100 0.100 ;
  LAYER metal2 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  LAYER metal3 ;
    RECT -0.300 -0.300 0.300 0.300 ;
END VIA2_1

VIA VIA3_1 DEFAULT
  LAYER via3 ;
    RECT -0.100 -0.100 0.100 0.100 ;
  LAYER metal3 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  LAYER topmetal ;
    RECT -0.300 -0.300 0.300 0.300 ;
END VIA3_1
