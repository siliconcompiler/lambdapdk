// //#############################################################################
// //# Function: 4-Input XOR Gate                                                #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_xor4 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     input  b,
//     input  c,
//     input  d,
//     output z
// );
// 
//     assign z = a ^ b ^ c ^ d;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
module la_xor4 (
    a,
    b,
    c,
    d,
    z
);
  wire _0_;
  wire _1_;
  (* src = "generated" *)
  input a;
  wire a;
  (* src = "generated" *)
  input b;
  wire b;
  (* src = "generated" *)
  input c;
  wire c;
  (* src = "generated" *)
  input d;
  wire d;
  (* src = "generated" *)
  output z;
  wire z;
  XOR2_X2 _2_ (
      .A(c),
      .B(d),
      .Z(_0_)
  );
  XNOR2_X2 _3_ (
      .A (b),
      .B (a),
      .ZN(_1_)
  );
  XNOR2_X2 _4_ (
      .A (_0_),
      .B (_1_),
      .ZN(z)
  );
endmodule
