// //#############################################################################
// //# Function: And-Or (ao211) Gate                                             #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_ao211 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a0,
//     input  a1,
//     input  b0,
//     input  c0,
//     output z
// );
// 
//     assign z = (a0 & a1) | b0 | c0;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_ao211.v:10.1-22.10" *)
module la_ao211 (
    a0,
    a1,
    b0,
    c0,
    z
);
  wire _0_;
  (* src = "inputs/la_ao211.v:13.12-13.14" *)
  input a0;
  wire a0;
  (* src = "inputs/la_ao211.v:14.12-14.14" *)
  input a1;
  wire a1;
  (* src = "inputs/la_ao211.v:15.12-15.14" *)
  input b0;
  wire b0;
  (* src = "inputs/la_ao211.v:16.12-16.14" *)
  input c0;
  wire c0;
  (* src = "inputs/la_ao211.v:17.12-17.13" *)
  output z;
  wire z;
  AOI211_X2 _1_ (
      .A (b0),
      .B (c0),
      .C1(a1),
      .C2(a0),
      .ZN(_0_)
  );
  INV_X1 _2_ (
      .A (_0_),
      .ZN(z)
  );
endmodule
