// //#############################################################################
// //# Function: 3-Input XOR Gate                                                #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_xor3 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     input  b,
//     input  c,
//     output z
// );
// 
//   assign z = a ^ b ^ c;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_xor3.v:10.1-21.10" *)
module la_xor3 (
    a,
    b,
    c,
    z
);
  (* src = "inputs/la_xor3.v:13.12-13.13" *)
  input a;
  wire a;
  (* src = "inputs/la_xor3.v:14.12-14.13" *)
  input b;
  wire b;
  (* src = "inputs/la_xor3.v:15.12-15.13" *)
  input c;
  wire c;
  (* src = "inputs/la_xor3.v:16.12-16.13" *)
  output z;
  wire z;
  gf180mcu_fd_sc_mcu7t5v0__xor3_2 _0_ (
      .A1(b),
      .A2(a),
      .A3(c),
      .Z (z)
  );
endmodule
