// //#############################################################################
// //# Function: Carry Save Adder (4:2) (aka 5:3)                                #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_csa42 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     input  b,
//     input  c,
//     input  d,
//     input  cin,
//     output sum,
//     output carry,
//     output cout
// );
// 
//     assign cout   = (a & b) | (b & c) | (a & c);
//     assign sumint = a ^ b ^ c;
//     assign sum    = cin ^ d ^ sumint;
//     assign carry  = (cin & d) | (cin & sumint) | (d & sumint);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
module la_csa42 (
    a,
    b,
    c,
    d,
    cin,
    sum,
    carry,
    cout
);
  (* force_downto = 32'b00000000000000000000000000000001 *) (* src = "generated" *)
  wire _00_;
  (* force_downto = 32'b00000000000000000000000000000001 *) (* src = "generated" *)
  wire _01_;
  (* force_downto = 32'b00000000000000000000000000000001 *) (* src = "generated" *)
  wire _02_;
  (* force_downto = 32'b00000000000000000000000000000001 *) (* src = "generated" *)
  wire _03_;
  (* force_downto = 32'b00000000000000000000000000000001 *) (* src = "generated" *)
  wire _04_;
  (* force_downto = 32'b00000000000000000000000000000001 *) (* src = "generated" *)
  wire _05_;
  (* force_downto = 32'b00000000000000000000000000000001 *) (* src = "generated" *)
  wire _06_;
  (* force_downto = 32'b00000000000000000000000000000001 *) (* src = "generated" *)
  wire _07_;
  (* force_downto = 32'b00000000000000000000000000000001 *) (* src = "generated" *)
  wire _08_;
  (* force_downto = 32'b00000000000000000000000000000001 *) (* src = "generated" *)
  wire _09_;
  (* src = "generated" *)
  input a;
  wire a;
  (* src = "generated" *)
  input b;
  wire b;
  (* src = "generated" *)
  input c;
  wire c;
  (* src = "generated" *)
  output carry;
  wire carry;
  (* src = "generated" *)
  input cin;
  wire cin;
  (* src = "generated" *)
  output cout;
  wire cout;
  (* src = "generated" *)
  input d;
  wire d;
  (* src = "generated" *)
  output sum;
  wire sum;
  INV_X2 _10_ (
      .A (a),
      .ZN(_00_)
  );
  INV_X2 _11_ (
      .A (d),
      .ZN(_05_)
  );
  INV_X2 _12_ (
      .A (b),
      .ZN(_01_)
  );
  INV_X2 _13_ (
      .A (cin),
      .ZN(_06_)
  );
  INV_X2 _14_ (
      .A (c),
      .ZN(_02_)
  );
  INV_X2 _15_ (
      .A (_04_),
      .ZN(_07_)
  );
  INV_X2 _16_ (
      .A (_09_),
      .ZN(sum)
  );
  INV_X2 _17_ (
      .A (_03_),
      .ZN(cout)
  );
  INV_X2 _18_ (
      .A (_08_),
      .ZN(carry)
  );
  (* module_not_derived = 32'b00000000000000000000000000000001 *) (* src = "generated" *)
  FA_X1 _19_ (
      .A (_00_),
      .B (_01_),
      .CI(_02_),
      .CO(_03_),
      .S (_04_)
  );
  (* module_not_derived = 32'b00000000000000000000000000000001 *) (* src = "generated" *)
  FA_X1 _20_ (
      .A (_05_),
      .B (_06_),
      .CI(_07_),
      .CO(_08_),
      .S (_09_)
  );
endmodule
