// //#############################################################################
// //# Function: 3-Input XOR Gate                                                #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_xor3 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     input  b,
//     input  c,
//     output z
// );
// 
//     assign z = a ^ b ^ c;
// 
// endmodule

/* Generated by Yosys 0.40+33 (git sha1 cd1fb8b15, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_xor3(a, b, c, z);
  wire _0_;
  input a;
  wire a;
  input b;
  wire b;
  input c;
  wire c;
  output z;
  wire z;
  sg13g2_xnor2_1 _1_ (
    .A(a),
    .B(c),
    .Y(_0_)
  );
  sg13g2_xnor2_1 _2_ (
    .A(b),
    .B(_0_),
    .Y(z)
  );
endmodule
