// //#############################################################################
// //# Function: 3-Input one-hot mux                                             #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_dmux3 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  sel0,
//     input  sel1,
//     input  sel2,
//     input  in0,
//     input  in1,
//     input  in2,
//     output out
// );
// 
//     assign out = (sel0 & in0) | (sel1 & in1) | (sel2 & in2);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
module la_dmux3 (
    sel0,
    sel1,
    sel2,
    in0,
    in1,
    in2,
    out
);
  wire _0_;
  wire _1_;
  (* src = "generated" *)
  input in0;
  wire in0;
  (* src = "generated" *)
  input in1;
  wire in1;
  (* src = "generated" *)
  input in2;
  wire in2;
  (* src = "generated" *)
  output out;
  wire out;
  (* src = "generated" *)
  input sel0;
  wire sel0;
  (* src = "generated" *)
  input sel1;
  wire sel1;
  (* src = "generated" *)
  input sel2;
  wire sel2;
  sg13g2_nand2_1 _2_ (
      .A(in1),
      .B(sel1),
      .Y(_0_)
  );
  sg13g2_a22oi_1 _3_ (
      .A1(in2),
      .A2(sel2),
      .B1(in0),
      .B2(sel0),
      .Y (_1_)
  );
  sg13g2_nand2_1 _4_ (
      .A(_0_),
      .B(_1_),
      .Y(out)
  );
endmodule
