// //#############################################################################
// //# Function: 3 Input Nand Gate                                               #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_nand3 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     input  b,
//     input  c,
//     output z
// );
// 
//     assign z = ~(a & b & c);
// 
// endmodule

/* Generated by Yosys 0.40+33 (git sha1 cd1fb8b15, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_nand3(a, b, c, z);
  input a;
  wire a;
  input b;
  wire b;
  input c;
  wire c;
  output z;
  wire z;
  sg13g2_nand3_1 _0_ (
    .A(b),
    .B(a),
    .C(c),
    .Y(z)
  );
endmodule
