# Copyright 2024 ZeroASIC Corp
# 
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
# 
#      https://www.apache.org/licenses/LICENSE-2.0
# 
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO BUMP10
  CLASS BUMP COVER ;
  FOREIGN BUMP10 0.0 0.0 ;
  ORIGIN 5.0 5.0 ;
  SYMMETRY X Y ;
  SIZE 10.00 BY 10.00 ;
  PIN PAD
    DIRECTION INOUT ;
    PORT
      LAYER topmetal ;
        POLYGON 2 -5 -2 -5 -5 -2 -5 2 -2 5 2 5 5 2 5 -2 ;
    END
  END PAD
END BUMP10

MACRO BUMP45
  CLASS BUMP COVER ;
  FOREIGN BUMP10 0.0 0.0 ;
  ORIGIN 14.0 14.0 ;
  SYMMETRY X Y ;
  SIZE 28.00 BY 28.00 ;
  PIN PAD
    DIRECTION INOUT ;
    PORT
      LAYER topmetal ;
        POLYGON 6 -14 -6 -14 -14 -6 -14 6 -6 14 6 14 14 6 14 -6 ;
    END
  END PAD
END BUMP45
