// //#############################################################################
// //# Function: 3-Input Exclusive-Nor Gate                                      #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_xnor3 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     input  b,
//     input  c,
//     output z
// );
// 
//     assign z = ~(a ^ b ^ c);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_xnor3.v:10.1-21.10" *)
module la_xnor3 (
    a,
    b,
    c,
    z
);
  wire _0_;
  (* src = "inputs/la_xnor3.v:13.12-13.13" *)
  input a;
  wire a;
  (* src = "inputs/la_xnor3.v:14.12-14.13" *)
  input b;
  wire b;
  (* src = "inputs/la_xnor3.v:15.12-15.13" *)
  input c;
  wire c;
  (* src = "inputs/la_xnor3.v:16.12-16.13" *)
  output z;
  wire z;
  sg13g2_xor2_1 _1_ (
      .A(a),
      .B(c),
      .X(_0_)
  );
  sg13g2_xnor2_1 _2_ (
      .A(b),
      .B(_0_),
      .Y(z)
  );
endmodule
