// //#############################################################################
// //# Function: Non-inverting buffer with supplies                              #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_pwrbuf #(
//     parameter TARGET = "DEFAULT",  // "SIM"
//     parameter PROP   = "DEFAULT"
// ) (
//     input  vdd,
//     input  vss,
//     input  a,
//     output z
// );
// 
//     generate
//         if (TARGET == "SIM") assign z = ((vdd === 1'b1) && (vss === 1'b0)) ? a : 1'bX;
//         else assign z = a;
//     endgenerate
// 
// endmodule

/* Generated by Yosys 0.40 (git sha1 a1bb0255d, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_pwrbuf(vdd, vss, a, z);
  input a;
  wire a;
  input vdd;
  wire vdd;
  input vss;
  wire vss;
  output z;
  wire z;
  assign z = a;
endmodule
