// Source ../.sc/cache/ihp130-68eebafcd9b2f5e92c69d37a8d3d90eb266550f5/ihp-sg13g2/libs.ref/sg13g2_io/lef/sg13g2_io.lef

(* blackbox *)
module sg13g2_Corner (
    inout iovdd,
    inout iovss,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_Filler200 (
    inout iovdd,
    inout iovss,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_Filler400 (
    inout iovdd,
    inout iovss,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_Filler1000 (
    inout iovdd,
    inout iovss,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_Filler2000 (
    inout iovdd,
    inout iovss,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_Filler4000 (
    inout iovdd,
    inout iovss,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_Filler10000 (
    inout iovdd,
    inout iovss,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadIn (
    inout iovdd,
    inout iovss,
    inout p2c,
    inout pad,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadOut4mA (
    inout c2p,
    inout iovdd,
    inout iovss,
    inout pad,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadOut16mA (
    inout c2p,
    inout iovdd,
    inout iovss,
    inout pad,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadOut30mA (
    inout c2p,
    inout iovdd,
    inout iovss,
    inout pad,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadTriOut4mA (
    inout c2p,
    inout c2p_en,
    inout iovdd,
    inout iovss,
    inout pad,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadTriOut16mA (
    inout c2p,
    inout c2p_en,
    inout iovdd,
    inout iovss,
    inout pad,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadTriOut30mA (
    inout c2p,
    inout c2p_en,
    inout iovdd,
    inout iovss,
    inout pad,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadInOut4mA (
    inout c2p,
    inout c2p_en,
    inout iovdd,
    inout iovss,
    inout p2c,
    inout pad,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadInOut16mA (
    inout c2p,
    inout c2p_en,
    inout iovdd,
    inout iovss,
    inout p2c,
    inout pad,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadInOut30mA (
    inout c2p,
    inout c2p_en,
    inout iovdd,
    inout iovss,
    inout p2c,
    inout pad,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadAnalog (
    inout iovdd,
    inout iovss,
    inout pad,
    inout padres,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadIOVss (
    inout iovdd,
    inout iovss,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadIOVdd (
    inout iovdd,
    inout iovss,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadVss (
    inout iovdd,
    inout iovss,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadVdd (
    inout iovdd,
    inout iovss,
    inout vdd,
    inout vss
);
endmodule
