// //#############################################################################
// //# Function: Or-And (oa33) Gate                                              #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_oa33 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a0,
//     input  a1,
//     input  a2,
//     input  b0,
//     input  b1,
//     input  b2,
//     output z
// );
// 
//     assign z = (a0 | a1 | a2) & (b0 | b1 | b2);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
(* keep_hierarchy *)
module la_oa33 (
    a0,
    a1,
    a2,
    b0,
    b1,
    b2,
    z
);
  (* src = "generated" *)
  input a0;
  wire a0;
  (* src = "generated" *)
  input a1;
  wire a1;
  (* src = "generated" *)
  input a2;
  wire a2;
  (* src = "generated" *)
  input b0;
  wire b0;
  (* src = "generated" *)
  input b1;
  wire b1;
  (* src = "generated" *)
  input b2;
  wire b2;
  (* src = "generated" *)
  output z;
  wire z;
  OA33x2_ASAP7_75t_R _0_ (
      .A1(a1),
      .A2(a0),
      .A3(a2),
      .B1(b1),
      .B2(b0),
      .B3(b2),
      .Y (z)
  );
endmodule
