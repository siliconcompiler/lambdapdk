// //#############################################################################
// //# Function: Power isolation circuit                                         #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_isohi #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  iso,  // isolation signal
//     input  in,   // input
//     output out   // out = iso | in
// );
// 
//     assign out = iso | in;
// 
// endmodule

/* Generated by Yosys 0.40 (git sha1 a1bb0255d, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_isohi(iso, in, out);
  input in;
  wire in;
  input iso;
  wire iso;
  output out;
  wire out;
  OR2x2_ASAP7_75t_SL _0_ (
    .A(in),
    .B(iso),
    .Y(out)
  );
endmodule
