// //#############################################################################
// //# Function: 2 Input Or Gate                                                 #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_or2 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     input  b,
//     output z
// );
// 
//   assign z = a | b;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_or2.v:10.1-20.10" *)
module la_or2 (
    a,
    b,
    z
);
  (* src = "inputs/la_or2.v:13.12-13.13" *)
  input a;
  wire a;
  (* src = "inputs/la_or2.v:14.12-14.13" *)
  input b;
  wire b;
  (* src = "inputs/la_or2.v:15.12-15.13" *)
  output z;
  wire z;
  OR2x2_ASAP7_75t_L _0_ (
      .A(b),
      .B(a),
      .Y(z)
  );
endmodule
