//#############################################################################
//# Function: Charge Keeper Cell                                              #
//# Copyright: Lambda Project Authors. All rights Reserved.                   #
//# License:  MIT (see LICENSE file in Lambda repository)                     #
//#############################################################################

module la_keeper #(
    parameter PROP = "DEFAULT"
) (
    inout z
);

endmodule
