// //#############################################################################
// //# Function: Carry Save Adder (4:2) (aka 5:3)                                #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_csa42 #(parameter PROP = "DEFAULT")  ( input  a,
//     input  b,
//     input  c,
//     input  d,
//     input  cin,
//     output sum,
//     output carry,
//     output cout
//     );
// 
//    assign cout   = (a & b) | (b & c) | (a & c);
//    assign sumint = a ^ b ^ c;
//    assign sum    = cin ^ d ^ sumint;
//    assign carry  = (cin & d) | (cin & sumint) | (d & sumint);
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_csa42(a, b, c, d, cin, sum, carry, cout);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  input a;
  wire a;
  input b;
  wire b;
  input c;
  wire c;
  output carry;
  wire carry;
  input cin;
  wire cin;
  output cout;
  wire cout;
  input d;
  wire d;
  output sum;
  wire sum;
  gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _10_ (
    .I(a),
    .ZN(_00_)
  );
  gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _11_ (
    .I(d),
    .ZN(_05_)
  );
  gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _12_ (
    .I(b),
    .ZN(_01_)
  );
  gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _13_ (
    .I(cin),
    .ZN(_06_)
  );
  gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _14_ (
    .I(c),
    .ZN(_02_)
  );
  gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _15_ (
    .I(_04_),
    .ZN(_07_)
  );
  gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _16_ (
    .I(_09_),
    .ZN(sum)
  );
  gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _17_ (
    .I(_03_),
    .ZN(cout)
  );
  gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _18_ (
    .I(_08_),
    .ZN(carry)
  );
  gf180mcu_fd_sc_mcu7t5v0__addf_1 _19_ (
    .A(_00_),
    .B(_01_),
    .CI(_02_),
    .CO(_03_),
    .S(_04_)
  );
  gf180mcu_fd_sc_mcu7t5v0__addf_1 _20_ (
    .A(_05_),
    .B(_06_),
    .CI(_07_),
    .CO(_08_),
    .S(_09_)
  );
endmodule
