// //#############################################################################
// //# Function:  Positive edge-triggered static D-type flop-flop with async     #
// //#            active low preset and scan input.                              #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_sdffsq #(parameter PROP = "DEFAULT")   (
//     input      d,
//     input      si,
//     input      se,
//     input      clk,
//     input      nset,
//     output reg q
//     );
// 
//    always @ (posedge clk or negedge nset)
//      if(!nset)
//        q <= 1'b1;
//      else
//        q <= se ? si : d;
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_sdffsq(d, si, se, clk, nset, q);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  input clk;
  wire clk;
  input d;
  wire d;
  input nset;
  wire nset;
  output q;
  wire q;
  input se;
  wire se;
  input si;
  wire si;
  INVx2_ASAP7_75t_L _06_ (
    .A(se),
    .Y(_04_)
  );
  AND2x4_ASAP7_75t_L _07_ (
    .A(si),
    .B(se),
    .Y(_03_)
  );
  AO21x1_ASAP7_75t_L _08_ (
    .A1(d),
    .A2(_04_),
    .B(_03_),
    .Y(_00_)
  );
  INVx2_ASAP7_75t_L _09_ (
    .A(nset),
    .Y(_02_)
  );
  INVx2_ASAP7_75t_L _10_ (
    .A(_01_),
    .Y(q)
  );
  ASYNC_DFFHx1_ASAP7_75t_L _11_ (
    .CLK(clk),
    .D(_00_),
    .QN(_01_),
    .RESET(_05_),
    .SET(_02_)
  );
  TIELOx1_ASAP7_75t_L _12_ (
    .L(_05_)
  );
endmodule
