// //#############################################################################
// //# Function: Dual data rate input buffer                                     #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_iddr #(parameter PROP = "DEFAULT")   (
//     input      clk,     // clock
//     input      in,      // data input sampled on both edges of clock
//     output reg outrise, // rising edge sample
//     output reg outfall  // falling edge sample
//     );
// 
//    // Negedge Sample
//    always @ (negedge clk)
//      outfall <= in;
// 
//    // Posedge Sample
//    reg 	       inrise;
//    always @ (posedge clk)
//      inrise <= in;
// 
//    // Posedge Latch (for hold)
//    always @ (clk or inrise)
//      if(~clk)
//        outrise <= inrise;
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_iddr(clk, in, outrise, outfall);
  wire _0_;
  input clk;
  wire clk;
  input in;
  wire in;
  wire inrise;
  output outfall;
  wire outfall;
  output outrise;
  wire outrise;
  sky130_fd_sc_hdll__inv_1 _1_ (
    .A(clk),
    .Y(_0_)
  );
  sky130_fd_sc_hdll__dlxtn_1 _2_ (
    .D(inrise),
    .GATE_N(clk),
    .Q(outrise)
  );
  sky130_fd_sc_hdll__dfxtp_1 _3_ (
    .CLK(clk),
    .D(in),
    .Q(inrise)
  );
  sky130_fd_sc_hdll__dfxtp_1 _4_ (
    .CLK(_0_),
    .D(in),
    .Q(outfall)
  );
endmodule
