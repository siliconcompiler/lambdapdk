// //#############################################################################
// //# Function: Carry Save Adder (4:2) (aka 5:3)                                #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_csa42 #(parameter PROP = "DEFAULT")  ( input  a,
//     input  b,
//     input  c,
//     input  d,
//     input  cin,
//     output sum,
//     output carry,
//     output cout
//     );
// 
//    assign cout   = (a & b) | (b & c) | (a & c);
//    assign sumint = a ^ b ^ c;
//    assign sum    = cin ^ d ^ sumint;
//    assign carry  = (cin & d) | (cin & sumint) | (d & sumint);
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_csa42(a, b, c, d, cin, sum, carry, cout);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  input a;
  wire a;
  input b;
  wire b;
  input c;
  wire c;
  output carry;
  wire carry;
  input cin;
  wire cin;
  output cout;
  wire cout;
  input d;
  wire d;
  output sum;
  wire sum;
  sky130_fd_sc_hdll__inv_1 _10_ (
    .A(a),
    .Y(_00_)
  );
  sky130_fd_sc_hdll__inv_1 _11_ (
    .A(d),
    .Y(_05_)
  );
  sky130_fd_sc_hdll__inv_1 _12_ (
    .A(b),
    .Y(_01_)
  );
  sky130_fd_sc_hdll__inv_1 _13_ (
    .A(cin),
    .Y(_06_)
  );
  sky130_fd_sc_hdll__inv_1 _14_ (
    .A(c),
    .Y(_02_)
  );
  sky130_fd_sc_hdll__inv_1 _15_ (
    .A(_04_),
    .Y(_07_)
  );
  sky130_fd_sc_hdll__inv_1 _16_ (
    .A(_09_),
    .Y(sum)
  );
  sky130_fd_sc_hdll__inv_1 _17_ (
    .A(_03_),
    .Y(cout)
  );
  sky130_fd_sc_hdll__inv_1 _18_ (
    .A(_08_),
    .Y(carry)
  );
  sky130_fd_sc_hdll__fa_1 _19_ (
    .A(_00_),
    .B(_01_),
    .CIN(_02_),
    .COUT(_03_),
    .SUM(_04_)
  );
  sky130_fd_sc_hdll__fa_1 _20_ (
    .A(_05_),
    .B(_06_),
    .CIN(_07_),
    .COUT(_08_),
    .SUM(_09_)
  );
endmodule
