// //#############################################################################
// //# Function: Carry Save Adder (3:2)                                          #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_csa32 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     input  b,
//     input  c,
//     output sum,
//     output carry
// );
// 
//     assign sum   = a ^ b ^ c;
//     assign carry = (a & b) | (b & c) | (c & a);
// 
// endmodule

/* Generated by Yosys 0.40+33 (git sha1 cd1fb8b15, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_csa32(a, b, c, sum, carry);
  wire _0_;
  wire _1_;
  wire _2_;
  input a;
  wire a;
  input b;
  wire b;
  input c;
  wire c;
  output carry;
  wire carry;
  output sum;
  wire sum;
  sg13g2_xnor2_1 _3_ (
    .A(b),
    .B(c),
    .Y(_0_)
  );
  sg13g2_xnor2_1 _4_ (
    .A(a),
    .B(_0_),
    .Y(sum)
  );
  sg13g2_nand2_1 _5_ (
    .A(b),
    .B(c),
    .Y(_1_)
  );
  sg13g2_o21ai_1 _6_ (
    .A1(b),
    .A2(c),
    .B1(a),
    .Y(_2_)
  );
  sg13g2_nand2_1 _7_ (
    .A(_1_),
    .B(_2_),
    .Y(carry)
  );
endmodule
