// //#############################################################################
// //# Function: Positive edge-triggered inverting static D-type flop-flop       #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_dffqn #(
//     parameter PROP = "DEFAULT"
// ) (
//     input d,
//     input clk,
//     output reg qn
// );
// 
//     always @(posedge clk) qn <= ~d;
// 
// endmodule

/* Generated by Yosys 0.40 (git sha1 a1bb0255d, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_dffqn(d, clk, qn);
  wire _0_;
  wire _1_;
  input clk;
  wire clk;
  input d;
  wire d;
  output qn;
  wire qn;
  INVx1_ASAP7_75t_R _2_ (
    .A(d),
    .Y(_0_)
  );
  INVx1_ASAP7_75t_R _3_ (
    .A(_1_),
    .Y(qn)
  );
  DFFHQNx1_ASAP7_75t_R _4_ (
    .CLK(clk),
    .D(_0_),
    .QN(_1_)
  );
endmodule
