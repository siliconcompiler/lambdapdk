// //#############################################################################
// //# Function: 7-Input one-hot mux                                             #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_dmux7 #(
//     parameter PROP = "DEFAULT"  // cell property
// ) (
//     input  sel6,
//     input  sel5,
//     input  sel4,
//     input  sel3,
//     input  sel2,
//     input  sel1,
//     input  sel0,
//     input  in6,
//     input  in5,
//     input  in4,
//     input  in3,
//     input  in2,
//     input  in1,
//     input  in0,
//     output out
// );
// 
//   assign out = (sel0 & in0) |
//         (sel1 & in1) |
//         (sel2 & in2) |
//         (sel3 & in3) |
//         (sel4 & in4) |
//         (sel5 & in5) |
//         (sel6 & in6);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_dmux7.v:10.1-38.10" *)
module la_dmux7 (
    sel6,
    sel5,
    sel4,
    sel3,
    sel2,
    sel1,
    sel0,
    in6,
    in5,
    in4,
    in3,
    in2,
    in1,
    in0,
    out
);
  wire _0_;
  wire _1_;
  wire _2_;
  (* src = "inputs/la_dmux7.v:26.12-26.15" *)
  input in0;
  wire in0;
  (* src = "inputs/la_dmux7.v:25.12-25.15" *)
  input in1;
  wire in1;
  (* src = "inputs/la_dmux7.v:24.12-24.15" *)
  input in2;
  wire in2;
  (* src = "inputs/la_dmux7.v:23.12-23.15" *)
  input in3;
  wire in3;
  (* src = "inputs/la_dmux7.v:22.12-22.15" *)
  input in4;
  wire in4;
  (* src = "inputs/la_dmux7.v:21.12-21.15" *)
  input in5;
  wire in5;
  (* src = "inputs/la_dmux7.v:20.12-20.15" *)
  input in6;
  wire in6;
  (* src = "inputs/la_dmux7.v:27.12-27.15" *)
  output out;
  wire out;
  (* src = "inputs/la_dmux7.v:19.12-19.16" *)
  input sel0;
  wire sel0;
  (* src = "inputs/la_dmux7.v:18.12-18.16" *)
  input sel1;
  wire sel1;
  (* src = "inputs/la_dmux7.v:17.12-17.16" *)
  input sel2;
  wire sel2;
  (* src = "inputs/la_dmux7.v:16.12-16.16" *)
  input sel3;
  wire sel3;
  (* src = "inputs/la_dmux7.v:15.12-15.16" *)
  input sel4;
  wire sel4;
  (* src = "inputs/la_dmux7.v:14.12-14.16" *)
  input sel5;
  wire sel5;
  (* src = "inputs/la_dmux7.v:13.12-13.16" *)
  input sel6;
  wire sel6;
  sky130_fd_sc_hd__a22oi_1 _3_ (
      .A1(in0),
      .A2(sel0),
      .B1(in3),
      .B2(sel3),
      .Y (_0_)
  );
  sky130_fd_sc_hd__a222oi_1 _4_ (
      .A1(in1),
      .A2(sel1),
      .B1(in2),
      .B2(sel2),
      .C1(in4),
      .C2(sel4),
      .Y (_1_)
  );
  sky130_fd_sc_hd__a22oi_1 _5_ (
      .A1(in5),
      .A2(sel5),
      .B1(in6),
      .B2(sel6),
      .Y (_2_)
  );
  sky130_fd_sc_hd__nand3_1 _6_ (
      .A(_0_),
      .B(_1_),
      .C(_2_),
      .Y(out)
  );
endmodule
