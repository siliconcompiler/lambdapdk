// //#############################################################################
// //# Function: 2-Input Inverting Mux                                           #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_muxi2 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  d0,
//     input  d1,
//     input  s,
//     output z
// );
// 
//     assign z = ~((d0 & ~s) | (d1 & s));
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_muxi2.v:10.1-21.10" *)
module la_muxi2 (
    d0,
    d1,
    s,
    z
);
  (* src = "inputs/la_muxi2.v:13.12-13.14" *)
  input d0;
  wire d0;
  (* src = "inputs/la_muxi2.v:14.12-14.14" *)
  input d1;
  wire d1;
  (* src = "inputs/la_muxi2.v:15.12-15.13" *)
  input s;
  wire s;
  (* src = "inputs/la_muxi2.v:16.12-16.13" *)
  output z;
  wire z;
  sky130_fd_sc_hdll__mux2i_2 _0_ (
      .A0(d0),
      .A1(d1),
      .S (s),
      .Y (z)
  );
endmodule
