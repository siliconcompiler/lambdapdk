// //#############################################################################
// //# Function: Carry Save Adder (4:2) (aka 5:3)                                #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_csa42 #(parameter PROP = "DEFAULT")  ( input  a,
//     input  b,
//     input  c,
//     input  d,
//     input  cin,
//     output sum,
//     output carry,
//     output cout
//     );
// 
//    assign cout   = (a & b) | (b & c) | (a & c);
//    assign sumint = a ^ b ^ c;
//    assign sum    = cin ^ d ^ sumint;
//    assign carry  = (cin & d) | (cin & sumint) | (d & sumint);
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_csa42(a, b, c, d, cin, sum, carry, cout);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  input a;
  wire a;
  input b;
  wire b;
  input c;
  wire c;
  output carry;
  wire carry;
  input cin;
  wire cin;
  output cout;
  wire cout;
  input d;
  wire d;
  output sum;
  wire sum;
  INVx2_ASAP7_75t_R _06_ (
    .A(a),
    .Y(_00_)
  );
  INVx2_ASAP7_75t_R _07_ (
    .A(d),
    .Y(_03_)
  );
  INVx2_ASAP7_75t_R _08_ (
    .A(b),
    .Y(_01_)
  );
  INVx2_ASAP7_75t_R _09_ (
    .A(cin),
    .Y(_04_)
  );
  INVx2_ASAP7_75t_R _10_ (
    .A(c),
    .Y(_02_)
  );
  FAx1_ASAP7_75t_R _11_ (
    .A(_00_),
    .B(_01_),
    .CI(_02_),
    .CON(cout),
    .SN(_05_)
  );
  FAx1_ASAP7_75t_R _12_ (
    .A(_03_),
    .B(_04_),
    .CI(_05_),
    .CON(carry),
    .SN(sum)
  );
endmodule
