// //#############################################################################
// //# Function: Or-And-Inverter (oai33) Gate                                    #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_oai33 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a0,
//     input  a1,
//     input  a2,
//     input  b0,
//     input  b1,
//     input  b2,
//     output z
// );
// 
//     assign z = ~((a0 | a1 | a2) & (b0 | b1 | b2));
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
(* keep_hierarchy *)
module la_oai33 (
    a0,
    a1,
    a2,
    b0,
    b1,
    b2,
    z
);
  wire _0_;
  (* src = "generated" *)
  input a0;
  wire a0;
  (* src = "generated" *)
  input a1;
  wire a1;
  (* src = "generated" *)
  input a2;
  wire a2;
  (* src = "generated" *)
  input b0;
  wire b0;
  (* src = "generated" *)
  input b1;
  wire b1;
  (* src = "generated" *)
  input b2;
  wire b2;
  (* src = "generated" *)
  output z;
  wire z;
  OA33x2_ASAP7_75t_L _1_ (
      .A1(b1),
      .A2(b0),
      .A3(b2),
      .B1(a1),
      .B2(a0),
      .B3(a2),
      .Y (_0_)
  );
  INVx2_ASAP7_75t_L _2_ (
      .A(_0_),
      .Y(z)
  );
endmodule
