// //#############################################################################
// //# Function:  Positive edge-triggered static D-type flop-flop with async     #
// //#            active low reset.                                              #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_dffrq #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      clk,
//     input      nreset,
//     output reg q
// );
// 
//     always @(posedge clk or negedge nreset)
//         if (!nreset) q <= 1'b0;
//         else q <= d;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
(* keep_hierarchy *)
module la_dffrq (
    d,
    clk,
    nreset,
    q
);
  (* unused_bits = "0" *)
  wire _0_;
  (* src = "generated" *)
  input clk;
  wire clk;
  (* src = "generated" *)
  input d;
  wire d;
  (* src = "generated" *)
  input nreset;
  wire nreset;
  (* src = "generated" *)
  output q;
  wire q;
  (* src = "generated" *)
  sg13g2_dfrbp_1 _1_ (
      .CLK(clk),
      .D(d),
      .Q(q),
      .Q_N(_0_),
      .RESET_B(nreset)
  );
endmodule
