// //#############################################################################
// //# Function: 2-Input Inverting Mux                                           #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_muxi2 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  d0,
//     input  d1,
//     input  s,
//     output z
// );
// 
//     assign z = ~((d0 & ~s) | (d1 & s));
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
(* keep_hierarchy *)
module la_muxi2 (
    d0,
    d1,
    s,
    z
);
  wire _0_;
  wire _1_;
  (* src = "generated" *)
  input d0;
  wire d0;
  (* src = "generated" *)
  input d1;
  wire d1;
  (* src = "generated" *)
  input s;
  wire s;
  (* src = "generated" *)
  output z;
  wire z;
  INVx1_ASAP7_75t_L _2_ (
      .A(d1),
      .Y(_0_)
  );
  NOR2x1_ASAP7_75t_L _3_ (
      .A(d0),
      .B(s),
      .Y(_1_)
  );
  AO21x1_ASAP7_75t_L _4_ (
      .A1(_0_),
      .A2(s),
      .B (_1_),
      .Y (z)
  );
endmodule
