// //#############################################################################
// //# Function: Positive edge-triggered inverting static D-type flop-flop       #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_dffqn #(parameter PROP = "DEFAULT")   (
//     input  	d,
//     input  	clk,
//     output reg  qn
//     );
// 
//    always @ (posedge clk)
//      qn <= ~d;
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_dffqn(d, clk, qn);
  wire _0_;
  input clk;
  wire clk;
  input d;
  wire d;
  output qn;
  wire qn;
  sky130_fd_sc_hdll__inv_1 _1_ (
    .A(d),
    .Y(_0_)
  );
  sky130_fd_sc_hdll__dfxtp_1 _2_ (
    .CLK(clk),
    .D(_0_),
    .Q(qn)
  );
endmodule
