// //#############################################################################
// //# Function: Synchronizer with async reset                                   #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// module la_drsync
//   #(parameter PROP = "DEFAULT")
//    (
//     input  clk,    // clock
//     input  in,     // input data
//     input  nreset, // async active low reset
//     output out     // synchronized data
//     );
// 
//    localparam STAGES=2;
// 
//    reg [STAGES-1:0] shiftreg;
// 
//    always @ (posedge clk or negedge nreset)
//      if(!nreset)
//        shiftreg[STAGES-1:0] <= 'b0;
//      else
//        shiftreg[STAGES-1:0] <= {shiftreg[STAGES-2:0],in};
// 
//    assign out = shiftreg[STAGES-1];
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_drsync(clk, in, nreset, out);
  input clk;
  wire clk;
  input in;
  wire in;
  input nreset;
  wire nreset;
  output out;
  wire out;
  wire \shiftreg[0] ;
  gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 _0_ (
    .CLK(clk),
    .D(in),
    .Q(\shiftreg[0] ),
    .RN(nreset)
  );
  gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 _1_ (
    .CLK(clk),
    .D(\shiftreg[0] ),
    .Q(out),
    .RN(nreset)
  );
endmodule
