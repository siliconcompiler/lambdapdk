//#############################################################################
//# Function: Antenna Diode                                                   #
//# Copyright: Lambda Project Authors. All rights Reserved.                   #
//# License:  MIT (see LICENSE file in Lambda repository)                     #
//#############################################################################

(* keep_hierarchy *)
module la_antenna #(
    parameter PROP = "DEFAULT"
) (
    input  vss,
    output z
);

  sky130_fd_sc_hd__diode_2 u0 (
      .DIODE(z),
      .VGND (vss)
  );

endmodule
