module $_DLATCH_P_(input E, input D, output Q);
    gf180mcu_fd_sc_mcu9t5v0__latq_1 _TECHMAP_REPLACE_ (
        .D(D),
        .E(E),
        .Q(Q)
        );
endmodule

module $_DLATCH_N_(input E, input D, output Q);
    gf180mcu_fd_sc_mcu9t5v0__latq_1 _TECHMAP_REPLACE_ (
        .D(D),
        .E(~E),
        .Q(Q)
        );
endmodule
