// //#############################################################################
// //# Function: 4-Input one-hot mux                                             #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_dmux4 #(
//     parameter PROP = "DEFAULT"  // cell property
// ) (
//     input  sel3,
//     input  sel2,
//     input  sel1,
//     input  sel0,
//     input  in3,
//     input  in2,
//     input  in1,
//     input  in0,
//     output out
// );
// 
//     assign out = (sel0 & in0) | (sel1 & in1) | (sel2 & in2) | (sel3 & in3);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
module la_dmux4 (
    sel3,
    sel2,
    sel1,
    sel0,
    in3,
    in2,
    in1,
    in0,
    out
);
  wire _0_;
  wire _1_;
  (* src = "generated" *)
  input in0;
  wire in0;
  (* src = "generated" *)
  input in1;
  wire in1;
  (* src = "generated" *)
  input in2;
  wire in2;
  (* src = "generated" *)
  input in3;
  wire in3;
  (* src = "generated" *)
  output out;
  wire out;
  (* src = "generated" *)
  input sel0;
  wire sel0;
  (* src = "generated" *)
  input sel1;
  wire sel1;
  (* src = "generated" *)
  input sel2;
  wire sel2;
  (* src = "generated" *)
  input sel3;
  wire sel3;
  AOI22_X2 _2_ (
      .A1(in0),
      .A2(sel0),
      .B1(in2),
      .B2(sel2),
      .ZN(_0_)
  );
  AOI22_X2 _3_ (
      .A1(in1),
      .A2(sel1),
      .B1(in3),
      .B2(sel3),
      .ZN(_1_)
  );
  NAND2_X1 _4_ (
      .A1(_0_),
      .A2(_1_),
      .ZN(out)
  );
endmodule
