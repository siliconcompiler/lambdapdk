* NGSPICE file created from gf180mcu_fd_ip_sram__sram64x8m8wm1.ext - technology: gf180mcuA

.subckt nmos_5p0431058998329_64x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=0.96u l=0.6u
.ends

.subckt nmos_1p2$$46563372_64x8m81 nmos_5p0431058998329_64x8m81_0/S nmos_5p0431058998329_64x8m81_0/D
+ a_n31_n74# VSUBS
Xnmos_5p0431058998329_64x8m81_0 nmos_5p0431058998329_64x8m81_0/D a_n31_n74# nmos_5p0431058998329_64x8m81_0/S
+ VSUBS nmos_5p0431058998329_64x8m81
.ends

.subckt pmos_5p04310589983278_64x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=0.9u l=1.2u
.ends

.subckt nmos_5p04310589983298_64x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=0.6u l=1u
.ends

.subckt pmos_5p04310589983291_64x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=22.68u l=0.6u
.ends

.subckt pmos_1p2$$47815724_64x8m81 pmos_5p04310589983291_64x8m81_0/D w_n286_n141#
+ pmos_5p04310589983291_64x8m81_0/S a_n31_n74#
Xpmos_5p04310589983291_64x8m81_0 w_n286_n141# pmos_5p04310589983291_64x8m81_0/D a_n31_n74#
+ pmos_5p04310589983291_64x8m81_0/S pmos_5p04310589983291_64x8m81
.ends

.subckt pmos_5p04310589983287_64x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.89u l=0.6u
.ends

.subckt pmos_5p04310589983292_64x8m81 w_n208_n120# D a_2016_n44# a_0_n44# a_896_n44#
+ a_672_n44# S a_1792_n44# a_448_n44# a_224_n44# a_1568_n44# a_1344_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X5 S a_2016_n44# D w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X6 S a_1120_n44# D w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X7 D a_1344_n44# S w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X8 S a_1568_n44# D w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X9 D a_1792_n44# S w_n208_n120# pmos_6p0 w=12.48u l=0.6u
.ends

.subckt nmos_5p04310589983293_64x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=0.6u l=1.2u
.ends

.subckt pmos_5p04310589983296_64x8m81 a_2464_n44# w_n208_n120# D a_2240_n44# a_3584_n44#
+ a_2016_n44# a_3360_n44# a_3136_n44# a_2912_n44# a_0_n44# a_4256_n44# a_4032_n44#
+ a_3808_n44# a_896_n44# a_672_n44# S a_1792_n44# a_448_n44# a_224_n44# a_1568_n44#
+ a_1344_n44# a_1120_n44# a_2688_n44#
X0 D a_4032_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X1 S a_4256_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X2 S a_224_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X3 D a_448_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X4 D a_0_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X5 S a_2912_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X6 D a_3136_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X7 S a_672_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X8 D a_896_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X9 S a_3360_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X10 S a_2016_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X11 D a_3584_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X12 D a_2240_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X13 S a_2464_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X14 D a_2688_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X15 S a_1120_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X16 D a_1344_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X17 S a_1568_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X18 D a_1792_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X19 S a_3808_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
.ends

.subckt nmos_5p04310589983297_64x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=0.75u l=0.6u
.ends

.subckt pmos_5p0431058998323_64x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=1.14u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.14u l=0.6u
.ends

.subckt pmos_1p2$$46273580_64x8m81 pmos_5p0431058998323_64x8m81_0/D a_193_n74# w_n286_n142#
+ pmos_5p0431058998323_64x8m81_0/S a_n31_n74#
Xpmos_5p0431058998323_64x8m81_0 w_n286_n142# pmos_5p0431058998323_64x8m81_0/D a_n31_n74#
+ pmos_5p0431058998323_64x8m81_0/S a_193_n74# pmos_5p0431058998323_64x8m81
.ends

.subckt nmos_5p0431058998325_64x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
.ends

.subckt nmos_1p2$$46551084_64x8m81 nmos_5p0431058998325_64x8m81_0/D a_n31_n73# nmos_5p0431058998325_64x8m81_0/S
+ VSUBS
Xnmos_5p0431058998325_64x8m81_0 nmos_5p0431058998325_64x8m81_0/D a_n31_n73# nmos_5p0431058998325_64x8m81_0/S
+ VSUBS nmos_5p0431058998325_64x8m81
.ends

.subckt pmos_5p04310589983241_64x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=0.96u l=0.6u
.ends

.subckt nmos_5p04310589983279_64x8m81 D a_2016_n44# a_0_n44# a_896_n44# a_672_n44#
+ S a_1792_n44# a_448_n44# a_224_n44# a_1568_n44# a_1344_n44# a_1120_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=1.92u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=1.92u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=1.92u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=1.92u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=1.92u l=0.6u
X5 S a_2016_n44# D VSUBS nmos_6p0 w=1.92u l=0.6u
X6 S a_1120_n44# D VSUBS nmos_6p0 w=1.92u l=0.6u
X7 D a_1344_n44# S VSUBS nmos_6p0 w=1.92u l=0.6u
X8 S a_1568_n44# D VSUBS nmos_6p0 w=1.92u l=0.6u
X9 D a_1792_n44# S VSUBS nmos_6p0 w=1.92u l=0.6u
.ends

.subckt pmos_5p04310589983214_64x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
.ends

.subckt pmos_1p2$$202586156_64x8m81 pmos_5p04310589983214_64x8m81_0/S w_n286_n141#
+ pmos_5p04310589983214_64x8m81_0/D a_n31_n74#
Xpmos_5p04310589983214_64x8m81_0 w_n286_n141# pmos_5p04310589983214_64x8m81_0/D a_n31_n74#
+ pmos_5p04310589983214_64x8m81_0/S pmos_5p04310589983214_64x8m81
.ends

.subckt nmos_5p04310589983280_64x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=1.2u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=1.2u l=0.6u
.ends

.subckt pmos_5p04310589983283_64x8m81 w_n208_n120# D a_0_n44# a_896_n44# a_672_n44#
+ S a_448_n44# a_224_n44# a_1344_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.2u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=2.2u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.2u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=2.2u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=2.2u l=0.6u
X5 S a_1120_n44# D w_n208_n120# pmos_6p0 w=2.2u l=0.6u
X6 D a_1344_n44# S w_n208_n120# pmos_6p0 w=2.2u l=0.6u
.ends

.subckt pmos_5p04310589983282_64x8m81 w_n208_n120# D a_0_n44# a_896_n44# a_672_n44#
+ S a_448_n44# a_224_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.48u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=2.48u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.48u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=2.48u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=2.48u l=0.6u
X5 S a_1120_n44# D w_n208_n120# pmos_6p0 w=2.48u l=0.6u
.ends

.subckt nmos_5p04310589983239_64x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
.ends

.subckt pmos_5p04310589983220_64x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
.ends

.subckt pmos_1p2$$202587180_64x8m81 pmos_5p04310589983214_64x8m81_0/S w_n286_n141#
+ pmos_5p04310589983214_64x8m81_0/D a_n31_n74#
Xpmos_5p04310589983214_64x8m81_0 w_n286_n141# pmos_5p04310589983214_64x8m81_0/D a_n31_n74#
+ pmos_5p04310589983214_64x8m81_0/S pmos_5p04310589983214_64x8m81
.ends

.subckt pmos_5p04310589983281_64x8m81 w_n208_n120# D a_2016_n44# a_0_n44# a_896_n44#
+ a_672_n44# S a_1792_n44# a_448_n44# a_224_n44# a_1568_n44# a_1344_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X5 S a_2016_n44# D w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X6 S a_1120_n44# D w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X7 D a_1344_n44# S w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X8 S a_1568_n44# D w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X9 D a_1792_n44# S w_n208_n120# pmos_6p0 w=4.72u l=0.6u
.ends

.subckt nmos_5p04310589983286_64x8m81 D a_0_n44# S a_448_n44# a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2u l=0.6u
.ends

.subckt pmos_5p04310589983284_64x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.84u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.84u l=0.6u
.ends

.subckt nmos_5p04310589983285_64x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# a_1344_n44# a_1120_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=0.89u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=0.89u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=0.89u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=0.89u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=0.89u l=0.6u
X5 S a_1120_n44# D VSUBS nmos_6p0 w=0.89u l=0.6u
X6 D a_1344_n44# S VSUBS nmos_6p0 w=0.89u l=0.6u
.ends

.subckt nmos_1p2$$202595372_64x8m81 nmos_5p0431058998329_64x8m81_0/S nmos_5p0431058998329_64x8m81_0/D
+ a_n31_n73# VSUBS
Xnmos_5p0431058998329_64x8m81_0 nmos_5p0431058998329_64x8m81_0/D a_n31_n73# nmos_5p0431058998329_64x8m81_0/S
+ VSUBS nmos_5p0431058998329_64x8m81
.ends

.subckt nmos_1p2$$202596396_64x8m81 nmos_5p0431058998329_64x8m81_0/S nmos_5p0431058998329_64x8m81_0/D
+ a_n31_n73# VSUBS
Xnmos_5p0431058998329_64x8m81_0 nmos_5p0431058998329_64x8m81_0/D a_n31_n73# nmos_5p0431058998329_64x8m81_0/S
+ VSUBS nmos_5p0431058998329_64x8m81
.ends

.subckt wen_v2_64x8m81 wen GWE clk vss IGWEN vdd nmos_5p0431058998329_64x8m81_4/D
Xpmos_5p04310589983241_64x8m81_1 vdd pmos_5p04310589983241_64x8m81_1/D nmos_5p0431058998329_64x8m81_3/D
+ nmos_5p0431058998325_64x8m81_0/D pmos_5p04310589983241_64x8m81
Xnmos_5p04310589983279_64x8m81_0 GWE pmos_5p04310589983283_64x8m81_0/D pmos_5p04310589983283_64x8m81_0/D
+ pmos_5p04310589983283_64x8m81_0/D pmos_5p04310589983283_64x8m81_0/D vss pmos_5p04310589983283_64x8m81_0/D
+ pmos_5p04310589983283_64x8m81_0/D pmos_5p04310589983283_64x8m81_0/D pmos_5p04310589983283_64x8m81_0/D
+ pmos_5p04310589983283_64x8m81_0/D pmos_5p04310589983283_64x8m81_0/D vss nmos_5p04310589983279_64x8m81
Xnmos_5p0431058998329_64x8m81_3 nmos_5p0431058998329_64x8m81_3/D clk vss vss nmos_5p0431058998329_64x8m81
Xnmos_5p0431058998329_64x8m81_4 nmos_5p0431058998329_64x8m81_4/D nmos_5p0431058998329_64x8m81_3/D
+ vss vss nmos_5p0431058998329_64x8m81
Xnmos_5p04310589983279_64x8m81_1 IGWEN pmos_5p04310589983282_64x8m81_0/D pmos_5p04310589983282_64x8m81_0/D
+ pmos_5p04310589983282_64x8m81_0/D pmos_5p04310589983282_64x8m81_0/D vss pmos_5p04310589983282_64x8m81_0/D
+ pmos_5p04310589983282_64x8m81_0/D pmos_5p04310589983282_64x8m81_0/D pmos_5p04310589983282_64x8m81_0/D
+ pmos_5p04310589983282_64x8m81_0/D pmos_5p04310589983282_64x8m81_0/D vss nmos_5p04310589983279_64x8m81
Xpmos_1p2$$202586156_64x8m81_0 pmos_5p04310589983241_64x8m81_1/D vdd vdd pmos_5p04310589983214_64x8m81_2/S
+ pmos_1p2$$202586156_64x8m81
Xnmos_5p04310589983280_64x8m81_0 pmos_5p04310589983284_64x8m81_0/D pmos_5p04310589983214_64x8m81_2/S
+ vss pmos_5p04310589983214_64x8m81_2/S vss nmos_5p04310589983280_64x8m81
Xpmos_5p04310589983283_64x8m81_0 vdd pmos_5p04310589983283_64x8m81_0/D nmos_5p0431058998329_64x8m81_1/S
+ nmos_5p0431058998329_64x8m81_1/S nmos_5p0431058998329_64x8m81_1/S vdd nmos_5p0431058998329_64x8m81_1/S
+ nmos_5p0431058998329_64x8m81_1/S nmos_5p0431058998329_64x8m81_1/S nmos_5p0431058998329_64x8m81_1/S
+ pmos_5p04310589983283_64x8m81
Xpmos_5p04310589983282_64x8m81_0 vdd pmos_5p04310589983282_64x8m81_0/D wen wen wen
+ vdd wen wen wen pmos_5p04310589983282_64x8m81
Xnmos_5p04310589983239_64x8m81_0 pmos_5p04310589983284_64x8m81_0/D nmos_5p0431058998329_64x8m81_4/D
+ nmos_5p0431058998329_64x8m81_1/S nmos_5p0431058998329_64x8m81_4/D vss nmos_5p04310589983239_64x8m81
Xpmos_5p04310589983220_64x8m81_0 vdd pmos_5p04310589983284_64x8m81_0/D nmos_5p0431058998329_64x8m81_3/D
+ nmos_5p0431058998329_64x8m81_1/S nmos_5p0431058998329_64x8m81_3/D pmos_5p04310589983220_64x8m81
Xpmos_1p2$$202587180_64x8m81_0 nmos_5p0431058998329_64x8m81_2/S vdd nmos_5p0431058998325_64x8m81_0/D
+ nmos_5p0431058998329_64x8m81_4/D pmos_1p2$$202587180_64x8m81
Xpmos_5p04310589983214_64x8m81_0 vdd vdd pmos_5p04310589983283_64x8m81_0/D nmos_5p0431058998329_64x8m81_1/D
+ pmos_5p04310589983214_64x8m81
Xpmos_5p04310589983214_64x8m81_1 vdd nmos_5p0431058998329_64x8m81_3/D clk vdd pmos_5p04310589983214_64x8m81
Xpmos_5p04310589983214_64x8m81_2 vdd vdd nmos_5p0431058998325_64x8m81_0/D pmos_5p04310589983214_64x8m81_2/S
+ pmos_5p04310589983214_64x8m81
Xpmos_5p04310589983214_64x8m81_3 vdd vdd wen nmos_5p0431058998329_64x8m81_2/S pmos_5p04310589983214_64x8m81
Xpmos_5p04310589983281_64x8m81_0 vdd GWE pmos_5p04310589983283_64x8m81_0/D pmos_5p04310589983283_64x8m81_0/D
+ pmos_5p04310589983283_64x8m81_0/D pmos_5p04310589983283_64x8m81_0/D vdd pmos_5p04310589983283_64x8m81_0/D
+ pmos_5p04310589983283_64x8m81_0/D pmos_5p04310589983283_64x8m81_0/D pmos_5p04310589983283_64x8m81_0/D
+ pmos_5p04310589983283_64x8m81_0/D pmos_5p04310589983283_64x8m81_0/D pmos_5p04310589983281_64x8m81
Xpmos_5p04310589983214_64x8m81_4 vdd nmos_5p0431058998329_64x8m81_4/D nmos_5p0431058998329_64x8m81_3/D
+ vdd pmos_5p04310589983214_64x8m81
Xpmos_5p04310589983281_64x8m81_1 vdd IGWEN pmos_5p04310589983282_64x8m81_0/D pmos_5p04310589983282_64x8m81_0/D
+ pmos_5p04310589983282_64x8m81_0/D pmos_5p04310589983282_64x8m81_0/D vdd pmos_5p04310589983282_64x8m81_0/D
+ pmos_5p04310589983282_64x8m81_0/D pmos_5p04310589983282_64x8m81_0/D pmos_5p04310589983282_64x8m81_0/D
+ pmos_5p04310589983282_64x8m81_0/D pmos_5p04310589983282_64x8m81_0/D pmos_5p04310589983281_64x8m81
Xnmos_5p04310589983286_64x8m81_0 pmos_5p04310589983282_64x8m81_0/D wen vss wen wen
+ vss nmos_5p04310589983286_64x8m81
Xpmos_5p04310589983284_64x8m81_0 vdd pmos_5p04310589983284_64x8m81_0/D pmos_5p04310589983214_64x8m81_2/S
+ vdd pmos_5p04310589983214_64x8m81_2/S pmos_5p04310589983284_64x8m81
Xnmos_5p0431058998325_64x8m81_0 nmos_5p0431058998325_64x8m81_0/D nmos_5p0431058998329_64x8m81_3/D
+ nmos_5p0431058998329_64x8m81_2/S vss nmos_5p0431058998325_64x8m81
Xnmos_5p04310589983285_64x8m81_0 pmos_5p04310589983283_64x8m81_0/D nmos_5p0431058998329_64x8m81_1/S
+ nmos_5p0431058998329_64x8m81_1/S nmos_5p0431058998329_64x8m81_1/S vss nmos_5p0431058998329_64x8m81_1/S
+ nmos_5p0431058998329_64x8m81_1/S nmos_5p0431058998329_64x8m81_1/S nmos_5p0431058998329_64x8m81_1/S
+ vss nmos_5p04310589983285_64x8m81
Xnmos_5p0431058998329_64x8m81_0 vss pmos_5p04310589983283_64x8m81_0/D nmos_5p0431058998329_64x8m81_1/D
+ vss nmos_5p0431058998329_64x8m81
Xnmos_1p2$$202595372_64x8m81_0 pmos_5p04310589983214_64x8m81_2/S vss nmos_5p0431058998325_64x8m81_0/D
+ vss nmos_1p2$$202595372_64x8m81
Xnmos_1p2$$202595372_64x8m81_1 nmos_5p0431058998325_64x8m81_0/D pmos_5p04310589983241_64x8m81_1/D
+ nmos_5p0431058998329_64x8m81_4/D vss nmos_1p2$$202595372_64x8m81
Xnmos_5p0431058998329_64x8m81_1 nmos_5p0431058998329_64x8m81_1/D nmos_5p0431058998329_64x8m81_3/D
+ nmos_5p0431058998329_64x8m81_1/S vss nmos_5p0431058998329_64x8m81
Xpmos_5p04310589983241_64x8m81_0 vdd nmos_5p0431058998329_64x8m81_1/D nmos_5p0431058998329_64x8m81_4/D
+ nmos_5p0431058998329_64x8m81_1/S pmos_5p04310589983241_64x8m81
Xnmos_5p0431058998329_64x8m81_2 vss wen nmos_5p0431058998329_64x8m81_2/S vss nmos_5p0431058998329_64x8m81
Xnmos_1p2$$202596396_64x8m81_0 pmos_5p04310589983241_64x8m81_1/D vss pmos_5p04310589983214_64x8m81_2/S
+ vss nmos_1p2$$202596396_64x8m81
.ends

.subckt pmos_5p04310589983295_64x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=0.9u l=1u
.ends

.subckt nmos_5p04310589983257_64x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=1.36u l=0.6u
.ends

.subckt nmos_1p2$$47342636_64x8m81 nmos_5p04310589983257_64x8m81_0/S nmos_5p04310589983257_64x8m81_0/D
+ a_n31_n73# VSUBS
Xnmos_5p04310589983257_64x8m81_0 nmos_5p04310589983257_64x8m81_0/D a_n31_n73# nmos_5p04310589983257_64x8m81_0/S
+ VSUBS nmos_5p04310589983257_64x8m81
.ends

.subckt pmos_1p2$$46285868_64x8m81 pmos_5p04310589983214_64x8m81_0/S w_n286_n142#
+ pmos_5p04310589983214_64x8m81_0/D a_n31_n73#
Xpmos_5p04310589983214_64x8m81_0 w_n286_n142# pmos_5p04310589983214_64x8m81_0/D a_n31_n73#
+ pmos_5p04310589983214_64x8m81_0/S pmos_5p04310589983214_64x8m81
.ends

.subckt pmos_1p2$$47330348_64x8m81 pmos_5p04310589983241_64x8m81_0/D a_n31_n73# w_n286_n141#
+ pmos_5p04310589983241_64x8m81_0/S
Xpmos_5p04310589983241_64x8m81_0 w_n286_n141# pmos_5p04310589983241_64x8m81_0/D a_n31_n73#
+ pmos_5p04310589983241_64x8m81_0/S pmos_5p04310589983241_64x8m81
.ends

.subckt nmos_5p04310589983289_64x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=9.98u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=9.98u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=9.98u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=9.98u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=9.98u l=0.6u
.ends

.subckt nmos_1p2$$48306220_64x8m81 nmos_5p04310589983289_64x8m81_0/D a_865_n74# a_641_n74#
+ a_417_n74# a_193_n74# nmos_5p04310589983289_64x8m81_0/S a_n31_n74# VSUBS
Xnmos_5p04310589983289_64x8m81_0 nmos_5p04310589983289_64x8m81_0/D a_n31_n74# a_865_n74#
+ a_641_n74# nmos_5p04310589983289_64x8m81_0/S a_417_n74# a_193_n74# VSUBS nmos_5p04310589983289_64x8m81
.ends

.subckt pmos_5p04310589983277_64x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=3.77u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=3.77u l=0.6u
.ends

.subckt pmos_1p2$$48623660_64x8m81 pmos_5p04310589983277_64x8m81_0/S a_193_n74# pmos_5p04310589983277_64x8m81_0/D
+ w_n286_n142# a_n31_n74#
Xpmos_5p04310589983277_64x8m81_0 w_n286_n142# pmos_5p04310589983277_64x8m81_0/D a_n31_n74#
+ pmos_5p04310589983277_64x8m81_0/S a_193_n74# pmos_5p04310589983277_64x8m81
.ends

.subckt pmos_5p04310589983294_64x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=19.5u l=0.6u
.ends

.subckt pmos_1p2$$48624684_64x8m81 pmos_5p04310589983294_64x8m81_0/D w_n286_n141#
+ pmos_5p04310589983294_64x8m81_0/S a_n31_n74#
Xpmos_5p04310589983294_64x8m81_0 w_n286_n141# pmos_5p04310589983294_64x8m81_0/D a_n31_n74#
+ pmos_5p04310589983294_64x8m81_0/S pmos_5p04310589983294_64x8m81
.ends

.subckt nmos_5p04310589983288_64x8m81 a_2464_n44# D a_2240_n44# a_3584_n44# a_2016_n44#
+ a_3360_n44# a_3136_n44# a_2912_n44# a_0_n44# a_4256_n44# a_4032_n44# a_3808_n44#
+ a_896_n44# a_672_n44# S a_1792_n44# a_448_n44# a_224_n44# a_1568_n44# a_1344_n44#
+ a_1120_n44# a_2688_n44# VSUBS
X0 S a_4256_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X1 S a_224_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X2 D a_448_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X3 D a_0_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X4 S a_2912_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X5 D a_3136_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X6 S a_672_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X7 D a_896_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X8 S a_3360_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X9 S a_2016_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X10 D a_3584_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X11 D a_2240_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X12 S a_2464_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X13 D a_2688_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X14 S a_1120_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X15 D a_1344_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X16 S a_1568_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X17 D a_1792_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X18 S a_3808_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X19 D a_4032_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
.ends

.subckt nmos_1p2$$48308268_64x8m81 nmos_5p04310589983288_64x8m81_0/a_4032_n44# nmos_5p04310589983288_64x8m81_0/a_3808_n44#
+ nmos_5p04310589983288_64x8m81_0/a_1792_n44# nmos_5p04310589983288_64x8m81_0/a_1568_n44#
+ nmos_5p04310589983288_64x8m81_0/a_1344_n44# nmos_5p04310589983288_64x8m81_0/a_1120_n44#
+ nmos_5p04310589983288_64x8m81_0/a_2688_n44# nmos_5p04310589983288_64x8m81_0/a_2464_n44#
+ nmos_5p04310589983288_64x8m81_0/a_2240_n44# nmos_5p04310589983288_64x8m81_0/a_896_n44#
+ nmos_5p04310589983288_64x8m81_0/S nmos_5p04310589983288_64x8m81_0/a_672_n44# nmos_5p04310589983288_64x8m81_0/a_3584_n44#
+ nmos_5p04310589983288_64x8m81_0/a_0_n44# nmos_5p04310589983288_64x8m81_0/a_2016_n44#
+ nmos_5p04310589983288_64x8m81_0/a_3360_n44# nmos_5p04310589983288_64x8m81_0/a_448_n44#
+ nmos_5p04310589983288_64x8m81_0/a_224_n44# nmos_5p04310589983288_64x8m81_0/a_3136_n44#
+ nmos_5p04310589983288_64x8m81_0/a_2912_n44# nmos_5p04310589983288_64x8m81_0/a_4256_n44#
+ VSUBS nmos_5p04310589983288_64x8m81_0/D
Xnmos_5p04310589983288_64x8m81_0 nmos_5p04310589983288_64x8m81_0/a_2464_n44# nmos_5p04310589983288_64x8m81_0/D
+ nmos_5p04310589983288_64x8m81_0/a_2240_n44# nmos_5p04310589983288_64x8m81_0/a_3584_n44#
+ nmos_5p04310589983288_64x8m81_0/a_2016_n44# nmos_5p04310589983288_64x8m81_0/a_3360_n44#
+ nmos_5p04310589983288_64x8m81_0/a_3136_n44# nmos_5p04310589983288_64x8m81_0/a_2912_n44#
+ nmos_5p04310589983288_64x8m81_0/a_0_n44# nmos_5p04310589983288_64x8m81_0/a_4256_n44#
+ nmos_5p04310589983288_64x8m81_0/a_4032_n44# nmos_5p04310589983288_64x8m81_0/a_3808_n44#
+ nmos_5p04310589983288_64x8m81_0/a_896_n44# nmos_5p04310589983288_64x8m81_0/a_672_n44#
+ nmos_5p04310589983288_64x8m81_0/S nmos_5p04310589983288_64x8m81_0/a_1792_n44# nmos_5p04310589983288_64x8m81_0/a_448_n44#
+ nmos_5p04310589983288_64x8m81_0/a_224_n44# nmos_5p04310589983288_64x8m81_0/a_1568_n44#
+ nmos_5p04310589983288_64x8m81_0/a_1344_n44# nmos_5p04310589983288_64x8m81_0/a_1120_n44#
+ nmos_5p04310589983288_64x8m81_0/a_2688_n44# VSUBS nmos_5p04310589983288_64x8m81
.ends

.subckt nmos_1p2$$48629804_64x8m81 nmos_5p04310589983239_64x8m81_0/D a_193_n73# a_n31_n73#
+ nmos_5p04310589983239_64x8m81_0/S VSUBS
Xnmos_5p04310589983239_64x8m81_0 nmos_5p04310589983239_64x8m81_0/D a_n31_n73# nmos_5p04310589983239_64x8m81_0/S
+ a_193_n73# VSUBS nmos_5p04310589983239_64x8m81
.ends

.subckt pmos_5p04310589983251_64x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=5.67u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=5.67u l=0.6u
.ends

.subckt nmos_5p04310589983290_64x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=3.02u l=0.6u
.ends

.subckt nmos_1p2$$48302124_64x8m81 a_n31_n74# nmos_5p04310589983290_64x8m81_0/S nmos_5p04310589983290_64x8m81_0/D
+ VSUBS
Xnmos_5p04310589983290_64x8m81_0 nmos_5p04310589983290_64x8m81_0/D a_n31_n74# nmos_5p04310589983290_64x8m81_0/S
+ VSUBS nmos_5p04310589983290_64x8m81
.ends

.subckt gen_512x8_64x8m81 WEN GWE tblhl cen clk wen_v2_64x8m81_0/IGWEN pmos_5p04310589983292_64x8m81_0/D
+ wen_v2_64x8m81_0/nmos_5p0431058998329_64x8m81_4/D men VSS VDD
Xnmos_1p2$$46563372_64x8m81_1 pmos_1p2$$46273580_64x8m81_0/pmos_5p0431058998323_64x8m81_0/D
+ VSS pmos_5p04310589983251_64x8m81_0/D VSS nmos_1p2$$46563372_64x8m81
Xpmos_5p04310589983278_64x8m81_0 VDD pmos_5p04310589983278_64x8m81_0/D clk VDD pmos_5p04310589983278_64x8m81
Xnmos_1p2$$46563372_64x8m81_2 nmos_1p2$$46563372_64x8m81_2/nmos_5p0431058998329_64x8m81_0/S
+ pmos_1p2$$46273580_64x8m81_0/pmos_5p0431058998323_64x8m81_0/D nmos_1p2$$46563372_64x8m81_0/nmos_5p0431058998329_64x8m81_0/D
+ VSS nmos_1p2$$46563372_64x8m81
Xpmos_5p04310589983278_64x8m81_1 VDD pmos_5p04310589983278_64x8m81_1/D pmos_5p04310589983278_64x8m81_0/D
+ VDD pmos_5p04310589983278_64x8m81
Xnmos_5p04310589983298_64x8m81_0 pmos_5p04310589983295_64x8m81_0/D pmos_5p04310589983278_64x8m81_1/D
+ VSS VSS nmos_5p04310589983298_64x8m81
Xpmos_1p2$$47815724_64x8m81_0 VDD VDD pmos_1p2$$47815724_64x8m81_3/pmos_5p04310589983291_64x8m81_0/S
+ tblhl pmos_1p2$$47815724_64x8m81
Xpmos_1p2$$47815724_64x8m81_1 pmos_1p2$$47815724_64x8m81_3/pmos_5p04310589983291_64x8m81_0/S
+ VDD VDD pmos_1p2$$47815724_64x8m81_7/pmos_5p04310589983291_64x8m81_0/S pmos_1p2$$47815724_64x8m81
Xpmos_5p04310589983287_64x8m81_0 VDD pmos_5p04310589983287_64x8m81_0/D pmos_5p04310589983295_64x8m81_0/D
+ VDD pmos_5p04310589983287_64x8m81
Xpmos_1p2$$47815724_64x8m81_2 pmos_1p2$$47815724_64x8m81_3/pmos_5p04310589983291_64x8m81_0/S
+ VDD VDD tblhl pmos_1p2$$47815724_64x8m81
Xpmos_1p2$$47815724_64x8m81_3 VDD VDD pmos_1p2$$47815724_64x8m81_3/pmos_5p04310589983291_64x8m81_0/S
+ pmos_1p2$$47815724_64x8m81_7/pmos_5p04310589983291_64x8m81_0/S pmos_1p2$$47815724_64x8m81
Xpmos_1p2$$47815724_64x8m81_4 pmos_1p2$$47815724_64x8m81_7/pmos_5p04310589983291_64x8m81_0/S
+ VDD VDD pmos_1p2$$47815724_64x8m81_3/pmos_5p04310589983291_64x8m81_0/S pmos_1p2$$47815724_64x8m81
Xpmos_1p2$$47815724_64x8m81_5 pmos_1p2$$47815724_64x8m81_7/pmos_5p04310589983291_64x8m81_0/S
+ VDD VDD pmos_1p2$$48624684_64x8m81_2/pmos_5p04310589983294_64x8m81_0/S pmos_1p2$$47815724_64x8m81
Xpmos_5p04310589983292_64x8m81_0 VDD pmos_5p04310589983292_64x8m81_0/D pmos_1p2$$47815724_64x8m81_7/pmos_5p04310589983291_64x8m81_0/S
+ pmos_1p2$$47815724_64x8m81_7/pmos_5p04310589983291_64x8m81_0/S pmos_1p2$$47815724_64x8m81_7/pmos_5p04310589983291_64x8m81_0/S
+ pmos_1p2$$47815724_64x8m81_7/pmos_5p04310589983291_64x8m81_0/S VDD pmos_1p2$$47815724_64x8m81_7/pmos_5p04310589983291_64x8m81_0/S
+ pmos_1p2$$47815724_64x8m81_7/pmos_5p04310589983291_64x8m81_0/S pmos_1p2$$47815724_64x8m81_7/pmos_5p04310589983291_64x8m81_0/S
+ pmos_1p2$$47815724_64x8m81_7/pmos_5p04310589983291_64x8m81_0/S pmos_1p2$$47815724_64x8m81_7/pmos_5p04310589983291_64x8m81_0/S
+ pmos_1p2$$47815724_64x8m81_7/pmos_5p04310589983291_64x8m81_0/S pmos_5p04310589983292_64x8m81
Xpmos_1p2$$47815724_64x8m81_6 VDD VDD pmos_1p2$$47815724_64x8m81_7/pmos_5p04310589983291_64x8m81_0/S
+ pmos_1p2$$47815724_64x8m81_3/pmos_5p04310589983291_64x8m81_0/S pmos_1p2$$47815724_64x8m81
Xnmos_5p04310589983293_64x8m81_0 pmos_5p04310589983278_64x8m81_0/D clk VSS VSS nmos_5p04310589983293_64x8m81
Xpmos_5p04310589983296_64x8m81_0 pmos_5p04310589983292_64x8m81_0/D VDD men pmos_5p04310589983292_64x8m81_0/D
+ pmos_5p04310589983292_64x8m81_0/D pmos_5p04310589983292_64x8m81_0/D pmos_5p04310589983292_64x8m81_0/D
+ pmos_5p04310589983292_64x8m81_0/D pmos_5p04310589983292_64x8m81_0/D pmos_5p04310589983292_64x8m81_0/D
+ pmos_5p04310589983292_64x8m81_0/D pmos_5p04310589983292_64x8m81_0/D pmos_5p04310589983292_64x8m81_0/D
+ pmos_5p04310589983292_64x8m81_0/D pmos_5p04310589983292_64x8m81_0/D VDD pmos_5p04310589983292_64x8m81_0/D
+ pmos_5p04310589983292_64x8m81_0/D pmos_5p04310589983292_64x8m81_0/D pmos_5p04310589983292_64x8m81_0/D
+ pmos_5p04310589983292_64x8m81_0/D pmos_5p04310589983292_64x8m81_0/D pmos_5p04310589983292_64x8m81_0/D
+ pmos_5p04310589983296_64x8m81
Xpmos_1p2$$47815724_64x8m81_7 VDD VDD pmos_1p2$$47815724_64x8m81_7/pmos_5p04310589983291_64x8m81_0/S
+ pmos_1p2$$48624684_64x8m81_2/pmos_5p04310589983294_64x8m81_0/S pmos_1p2$$47815724_64x8m81
Xnmos_5p04310589983297_64x8m81_0 pmos_5p04310589983287_64x8m81_0/D pmos_5p04310589983295_64x8m81_0/D
+ VSS VSS nmos_5p04310589983297_64x8m81
Xnmos_5p04310589983293_64x8m81_1 pmos_5p04310589983278_64x8m81_1/D pmos_5p04310589983278_64x8m81_0/D
+ VSS VSS nmos_5p04310589983293_64x8m81
Xpmos_1p2$$46273580_64x8m81_0 pmos_1p2$$46273580_64x8m81_0/pmos_5p0431058998323_64x8m81_0/D
+ pmos_5p04310589983251_64x8m81_0/D VDD VDD pmos_5p04310589983251_64x8m81_0/D pmos_1p2$$46273580_64x8m81
Xnmos_1p2$$46551084_64x8m81_0 cen nmos_1p2$$47342636_64x8m81_1/nmos_5p04310589983257_64x8m81_0/S
+ nmos_1p2$$46563372_64x8m81_2/nmos_5p0431058998329_64x8m81_0/S VSS nmos_1p2$$46551084_64x8m81
Xwen_v2_64x8m81_0 wen_v2_64x8m81_0/wen wen_v2_64x8m81_0/GWE clk VSS wen_v2_64x8m81_0/IGWEN
+ VDD wen_v2_64x8m81_0/nmos_5p0431058998329_64x8m81_4/D wen_v2_64x8m81
Xpmos_5p04310589983295_64x8m81_0 VDD pmos_5p04310589983295_64x8m81_0/D pmos_5p04310589983278_64x8m81_1/D
+ VDD pmos_5p04310589983295_64x8m81
Xnmos_1p2$$47342636_64x8m81_0 VSS nmos_1p2$$47342636_64x8m81_1/nmos_5p04310589983257_64x8m81_0/S
+ clk VSS nmos_1p2$$47342636_64x8m81
Xpmos_1p2$$46285868_64x8m81_0 VDD VDD nmos_1p2$$46563372_64x8m81_0/nmos_5p0431058998329_64x8m81_0/D
+ nmos_1p2$$47342636_64x8m81_1/nmos_5p04310589983257_64x8m81_0/S pmos_1p2$$46285868_64x8m81
Xnmos_1p2$$47342636_64x8m81_1 nmos_1p2$$47342636_64x8m81_1/nmos_5p04310589983257_64x8m81_0/S
+ VSS men VSS nmos_1p2$$47342636_64x8m81
Xpmos_1p2$$46285868_64x8m81_1 nmos_1p2$$46563372_64x8m81_2/nmos_5p0431058998329_64x8m81_0/S
+ VDD cen nmos_1p2$$46563372_64x8m81_0/nmos_5p0431058998329_64x8m81_0/D pmos_1p2$$46285868_64x8m81
Xpmos_1p2$$47330348_64x8m81_0 pmos_1p2$$46273580_64x8m81_0/pmos_5p0431058998323_64x8m81_0/D
+ nmos_1p2$$47342636_64x8m81_1/nmos_5p04310589983257_64x8m81_0/S VDD nmos_1p2$$46563372_64x8m81_2/nmos_5p0431058998329_64x8m81_0/S
+ pmos_1p2$$47330348_64x8m81
Xnmos_1p2$$48306220_64x8m81_0 pmos_5p04310589983292_64x8m81_0/D pmos_1p2$$47815724_64x8m81_7/pmos_5p04310589983291_64x8m81_0/S
+ pmos_1p2$$47815724_64x8m81_7/pmos_5p04310589983291_64x8m81_0/S pmos_1p2$$47815724_64x8m81_7/pmos_5p04310589983291_64x8m81_0/S
+ pmos_1p2$$47815724_64x8m81_7/pmos_5p04310589983291_64x8m81_0/S VSS pmos_1p2$$47815724_64x8m81_7/pmos_5p04310589983291_64x8m81_0/S
+ VSS nmos_1p2$$48306220_64x8m81
Xpmos_1p2$$48623660_64x8m81_0 VDD pmos_5p04310589983287_64x8m81_0/D pmos_1p2$$48623660_64x8m81_0/pmos_5p04310589983277_64x8m81_0/D
+ VDD pmos_5p04310589983287_64x8m81_0/D pmos_1p2$$48623660_64x8m81
Xpmos_1p2$$48624684_64x8m81_0 pmos_1p2$$48624684_64x8m81_2/pmos_5p04310589983294_64x8m81_0/S
+ VDD VDD pmos_5p04310589983251_64x8m81_0/D pmos_1p2$$48624684_64x8m81
Xnmos_1p2$$48308268_64x8m81_0 pmos_5p04310589983292_64x8m81_0/D pmos_5p04310589983292_64x8m81_0/D
+ pmos_5p04310589983292_64x8m81_0/D pmos_5p04310589983292_64x8m81_0/D pmos_5p04310589983292_64x8m81_0/D
+ pmos_5p04310589983292_64x8m81_0/D pmos_5p04310589983292_64x8m81_0/D pmos_5p04310589983292_64x8m81_0/D
+ pmos_5p04310589983292_64x8m81_0/D pmos_5p04310589983292_64x8m81_0/D VSS pmos_5p04310589983292_64x8m81_0/D
+ pmos_5p04310589983292_64x8m81_0/D pmos_5p04310589983292_64x8m81_0/D pmos_5p04310589983292_64x8m81_0/D
+ pmos_5p04310589983292_64x8m81_0/D pmos_5p04310589983292_64x8m81_0/D pmos_5p04310589983292_64x8m81_0/D
+ pmos_5p04310589983292_64x8m81_0/D pmos_5p04310589983292_64x8m81_0/D pmos_5p04310589983292_64x8m81_0/D
+ VSS men nmos_1p2$$48308268_64x8m81
Xpmos_1p2$$48624684_64x8m81_1 pmos_1p2$$48624684_64x8m81_2/pmos_5p04310589983294_64x8m81_0/S
+ VDD VDD pmos_1p2$$48623660_64x8m81_0/pmos_5p04310589983277_64x8m81_0/D pmos_1p2$$48624684_64x8m81
Xpmos_1p2$$48624684_64x8m81_2 VDD VDD pmos_1p2$$48624684_64x8m81_2/pmos_5p04310589983294_64x8m81_0/S
+ clk pmos_1p2$$48624684_64x8m81
Xnmos_1p2$$48629804_64x8m81_0 pmos_5p04310589983251_64x8m81_0/D nmos_1p2$$46563372_64x8m81_2/nmos_5p0431058998329_64x8m81_0/S
+ nmos_1p2$$46563372_64x8m81_2/nmos_5p0431058998329_64x8m81_0/S VSS VSS nmos_1p2$$48629804_64x8m81
Xpmos_5p04310589983251_64x8m81_0 VDD pmos_5p04310589983251_64x8m81_0/D nmos_1p2$$46563372_64x8m81_2/nmos_5p0431058998329_64x8m81_0/S
+ VDD nmos_1p2$$46563372_64x8m81_2/nmos_5p0431058998329_64x8m81_0/S pmos_5p04310589983251_64x8m81
Xnmos_1p2$$48302124_64x8m81_0 pmos_5p04310589983287_64x8m81_0/D VSS pmos_1p2$$48623660_64x8m81_0/pmos_5p04310589983277_64x8m81_0/D
+ VSS nmos_1p2$$48302124_64x8m81
Xnmos_1p2$$46563372_64x8m81_0 VSS nmos_1p2$$46563372_64x8m81_0/nmos_5p0431058998329_64x8m81_0/D
+ nmos_1p2$$47342636_64x8m81_1/nmos_5p04310589983257_64x8m81_0/S VSS nmos_1p2$$46563372_64x8m81
X0 VSS pmos_1p2$$47815724_64x8m81_3/pmos_5p04310589983291_64x8m81_0/S a_11293_484# VSS nmos_6p0 w=18.145u l=0.6u
X1 a_9646_262# pmos_1p2$$48623660_64x8m81_0/pmos_5p04310589983277_64x8m81_0/D VSS VSS nmos_6p0 w=22.68u l=0.6u
X2 pmos_1p2$$47815724_64x8m81_7/pmos_5p04310589983291_64x8m81_0/S pmos_1p2$$48624684_64x8m81_2/pmos_5p04310589983294_64x8m81_0/S a_10845_484# VSS nmos_6p0 w=18.145u l=0.6u
X3 a_12578_3205# tblhl pmos_1p2$$47815724_64x8m81_3/pmos_5p04310589983291_64x8m81_0/S VSS nmos_6p0 w=4.54u l=0.6u
X4 pmos_1p2$$48624684_64x8m81_2/pmos_5p04310589983294_64x8m81_0/S pmos_5p04310589983251_64x8m81_0/D a_9870_262# VSS nmos_6p0 w=22.68u l=0.6u
X5 a_11293_484# pmos_1p2$$48624684_64x8m81_2/pmos_5p04310589983294_64x8m81_0/S pmos_1p2$$47815724_64x8m81_7/pmos_5p04310589983291_64x8m81_0/S VSS nmos_6p0 w=18.145u l=0.6u
X6 a_12130_3205# pmos_1p2$$47815724_64x8m81_7/pmos_5p04310589983291_64x8m81_0/S VSS VSS nmos_6p0 w=4.54u l=0.6u
X7 a_10845_484# pmos_1p2$$47815724_64x8m81_3/pmos_5p04310589983291_64x8m81_0/S VSS VSS nmos_6p0 w=18.145u l=0.6u
X8 pmos_1p2$$47815724_64x8m81_3/pmos_5p04310589983291_64x8m81_0/S tblhl a_12130_3205# VSS nmos_6p0 w=4.54u l=0.6u
X9 nmos_1p2$$47342636_64x8m81_1/nmos_5p04310589983257_64x8m81_0/S clk a_5174_6131# VDD pmos_6p0 w=2.28u l=0.595u
X10 VSS pmos_1p2$$47815724_64x8m81_7/pmos_5p04310589983291_64x8m81_0/S a_12578_3205# VSS nmos_6p0 w=4.54u l=0.6u
X11 a_9870_262# clk a_9646_262# VSS nmos_6p0 w=22.68u l=0.6u
X12 a_5174_6131# men VDD VDD pmos_6p0 w=2.28u l=0.595u
.ends

.subckt pmos_5p0431058998324_64x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=13.61u l=0.6u
.ends

.subckt pmos_1p2$$46887980_64x8m81 pmos_5p0431058998324_64x8m81_0/D w_n286_n142# pmos_5p0431058998324_64x8m81_0/S
+ a_n31_n74#
Xpmos_5p0431058998324_64x8m81_0 w_n286_n142# pmos_5p0431058998324_64x8m81_0/D a_n31_n74#
+ pmos_5p0431058998324_64x8m81_0/S pmos_5p0431058998324_64x8m81
.ends

.subckt pmos_5p04310589983262_64x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=4.54u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=4.54u l=0.6u
.ends

.subckt pmos_1p2$$47331372_64x8m81 pmos_5p04310589983262_64x8m81_0/S a_n30_n74# w_n286_n142#
+ pmos_5p04310589983262_64x8m81_0/D a_194_n74#
Xpmos_5p04310589983262_64x8m81_0 w_n286_n142# pmos_5p04310589983262_64x8m81_0/D a_n30_n74#
+ pmos_5p04310589983262_64x8m81_0/S a_194_n74# pmos_5p04310589983262_64x8m81
.ends

.subckt pmos_1p2$$47330348_161_64x8m81 pmos_5p04310589983241_64x8m81_0/D a_n31_191#
+ w_n286_n141# pmos_5p04310589983241_64x8m81_0/S
Xpmos_5p04310589983241_64x8m81_0 w_n286_n141# pmos_5p04310589983241_64x8m81_0/D a_n31_191#
+ pmos_5p04310589983241_64x8m81_0/S pmos_5p04310589983241_64x8m81
.ends

.subckt nmos_1p2$$46551084_157_64x8m81 nmos_5p0431058998325_64x8m81_0/D a_n31_n74#
+ nmos_5p0431058998325_64x8m81_0/S VSUBS
Xnmos_5p0431058998325_64x8m81_0 nmos_5p0431058998325_64x8m81_0/D a_n31_n74# nmos_5p0431058998325_64x8m81_0/S
+ VSUBS nmos_5p0431058998325_64x8m81
.ends

.subckt nmos_5p04310589983263_64x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=1.82u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=1.82u l=0.6u
.ends

.subckt nmos_1p2$$47329324_64x8m81 a_194_n74# nmos_5p04310589983263_64x8m81_0/D nmos_5p04310589983263_64x8m81_0/S
+ a_n30_n74# VSUBS
Xnmos_5p04310589983263_64x8m81_0 nmos_5p04310589983263_64x8m81_0/D a_n30_n74# nmos_5p04310589983263_64x8m81_0/S
+ a_194_n74# VSUBS nmos_5p04310589983263_64x8m81
.ends

.subckt pmos_1p2$$46285868_160_64x8m81 pmos_5p04310589983214_64x8m81_0/S a_n31_n74#
+ w_n286_n142# pmos_5p04310589983214_64x8m81_0/D
Xpmos_5p04310589983214_64x8m81_0 w_n286_n142# pmos_5p04310589983214_64x8m81_0/D a_n31_n74#
+ pmos_5p04310589983214_64x8m81_0/S pmos_5p04310589983214_64x8m81
.ends

.subckt alatch_64x8m81 enb en ab a vss vdd
Xpmos_1p2$$47331372_64x8m81_0 vdd nmos_5p0431058998329_64x8m81_1/S vdd ab nmos_5p0431058998329_64x8m81_1/S
+ pmos_1p2$$47331372_64x8m81
Xpmos_1p2$$47330348_161_64x8m81_0 nmos_5p0431058998329_64x8m81_1/D en vdd nmos_5p0431058998329_64x8m81_1/S
+ pmos_1p2$$47330348_161_64x8m81
Xpmos_1p2$$47330348_161_64x8m81_1 vdd ab vdd nmos_5p0431058998329_64x8m81_1/D pmos_1p2$$47330348_161_64x8m81
Xnmos_1p2$$46551084_157_64x8m81_0 a en nmos_5p0431058998329_64x8m81_1/S vss nmos_1p2$$46551084_157_64x8m81
Xnmos_1p2$$47329324_64x8m81_0 nmos_5p0431058998329_64x8m81_1/S ab vss nmos_5p0431058998329_64x8m81_1/S
+ vss nmos_1p2$$47329324_64x8m81
Xpmos_1p2$$46285868_160_64x8m81_0 nmos_5p0431058998329_64x8m81_1/S enb vdd a pmos_1p2$$46285868_160_64x8m81
Xnmos_5p0431058998329_64x8m81_0 vss ab nmos_5p0431058998329_64x8m81_1/D vss nmos_5p0431058998329_64x8m81
Xnmos_5p0431058998329_64x8m81_1 nmos_5p0431058998329_64x8m81_1/D enb nmos_5p0431058998329_64x8m81_1/S
+ vss nmos_5p0431058998329_64x8m81
.ends

.subckt nmos_5p04310589983261_64x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=4.54u l=0.6u
.ends

.subckt nmos_1p2$$47514668_64x8m81 nmos_5p04310589983261_64x8m81_0/D a_n30_n73# nmos_5p04310589983261_64x8m81_0/S
+ VSUBS
Xnmos_5p04310589983261_64x8m81_0 nmos_5p04310589983261_64x8m81_0/D a_n30_n73# nmos_5p04310589983261_64x8m81_0/S
+ VSUBS nmos_5p04310589983261_64x8m81
.ends

.subckt ypredec1_bot_64x8m81 m1_n14_3279# m1_n14_2674# pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/S
+ alatch_64x8m81_0/vss m1_n14_2876# alatch_64x8m81_0/enb m1_n14_3078# m1_n14_3481#
+ alatch_64x8m81_0/vdd pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/D
+ m1_n14_2472# alatch_64x8m81_0/a pmos_1p2$$46887980_64x8m81_0/pmos_5p0431058998324_64x8m81_0/D
+ alatch_64x8m81_0/en
Xpmos_1p2$$46887980_64x8m81_0 pmos_1p2$$46887980_64x8m81_0/pmos_5p0431058998324_64x8m81_0/D
+ pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/S pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/S
+ pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/D pmos_1p2$$46887980_64x8m81
Xpmos_1p2$$46887980_64x8m81_1 pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/D
+ pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/S pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/S
+ alatch_64x8m81_0/ab pmos_1p2$$46887980_64x8m81
Xalatch_64x8m81_0 alatch_64x8m81_0/enb alatch_64x8m81_0/en alatch_64x8m81_0/ab alatch_64x8m81_0/a
+ alatch_64x8m81_0/vss alatch_64x8m81_0/vdd alatch_64x8m81
Xnmos_1p2$$47514668_64x8m81_0 pmos_1p2$$46887980_64x8m81_0/pmos_5p0431058998324_64x8m81_0/D
+ pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/D alatch_64x8m81_0/vss
+ alatch_64x8m81_0/vss nmos_1p2$$47514668_64x8m81
Xnmos_1p2$$47514668_64x8m81_1 pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/D
+ alatch_64x8m81_0/ab alatch_64x8m81_0/vss alatch_64x8m81_0/vss nmos_1p2$$47514668_64x8m81
.ends

.subckt nmos_5p04310589983260_64x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=1.91u l=0.6u
.ends

.subckt pmos_5p04310589983265_64x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=5.77u l=0.6u
.ends

.subckt pmos_1p2$$47820844_64x8m81 pmos_5p04310589983265_64x8m81_0/S w_n286_n141#
+ a_n30_n74# pmos_5p04310589983265_64x8m81_0/D
Xpmos_5p04310589983265_64x8m81_0 w_n286_n141# pmos_5p04310589983265_64x8m81_0/D a_n30_n74#
+ pmos_5p04310589983265_64x8m81_0/S pmos_5p04310589983265_64x8m81
.ends

.subckt pmos_5p04310589983264_64x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=5.67u l=0.6u
.ends

.subckt pmos_1p2$$47821868_64x8m81 pmos_5p04310589983264_64x8m81_0/S w_n286_n142#
+ pmos_5p04310589983264_64x8m81_0/D a_n31_n74#
Xpmos_5p04310589983264_64x8m81_0 w_n286_n142# pmos_5p04310589983264_64x8m81_0/D a_n31_n74#
+ pmos_5p04310589983264_64x8m81_0/S pmos_5p04310589983264_64x8m81
.ends

.subckt ypredec1_xa_64x8m81 m1_n58_n4290# m1_n58_n4895# m1_n58_n5097# m3_n1_n7124#
+ a_644_n6680# m1_n58_n4492# m1_n58_n4088# a_421_n4311# nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ a_n1_81# a_197_n5120# m1_n58_n4694# pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/S
+ M3_M2$$47819820_64x8m81_0/VSUBS
Xnmos_1p2$$46551084_64x8m81_1 M3_M2$$47819820_64x8m81_0/VSUBS pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/D
+ nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D M3_M2$$47819820_64x8m81_0/VSUBS
+ nmos_1p2$$46551084_64x8m81
Xnmos_1p2$$46551084_64x8m81_0 nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/D M3_M2$$47819820_64x8m81_0/VSUBS
+ M3_M2$$47819820_64x8m81_0/VSUBS nmos_1p2$$46551084_64x8m81
Xnmos_1p2$$46551084_64x8m81_2 nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/D M3_M2$$47819820_64x8m81_0/VSUBS
+ M3_M2$$47819820_64x8m81_0/VSUBS nmos_1p2$$46551084_64x8m81
Xpmos_1p2$$47820844_64x8m81_0 pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/S
+ pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/S pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/D
+ nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D pmos_1p2$$47820844_64x8m81
Xpmos_1p2$$47820844_64x8m81_1 pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/S
+ pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/S pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/D
+ nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D pmos_1p2$$47820844_64x8m81
Xpmos_1p2$$47821868_64x8m81_1 pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/D
+ pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/S pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/S
+ a_421_n4311# pmos_1p2$$47821868_64x8m81
Xpmos_1p2$$47821868_64x8m81_0 pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/S
+ pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/S pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/D
+ a_197_n5120# pmos_1p2$$47821868_64x8m81
Xpmos_1p2$$47820844_64x8m81_2 nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/S pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/D
+ pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/S pmos_1p2$$47820844_64x8m81
Xpmos_1p2$$47821868_64x8m81_2 pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/S
+ pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/S pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/D
+ a_644_n6680# pmos_1p2$$47821868_64x8m81
X0 pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/D a_644_n6680# a_542_n6607# M3_M2$$47819820_64x8m81_0/VSUBS nmos_3p3 w=6.81u l=0.6u
X1 a_318_n6607# a_197_n5120# M3_M2$$47819820_64x8m81_0/VSUBS M3_M2$$47819820_64x8m81_0/VSUBS nmos_3p3 w=6.81u l=0.6u
X2 a_542_n6607# a_421_n4311# a_318_n6607# M3_M2$$47819820_64x8m81_0/VSUBS nmos_3p3 w=6.81u l=0.6u
.ends

.subckt ypredec1_xax8_64x8m81 ypredec1_xa_64x8m81_1/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_xa_64x8m81_2/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ a_527_2758# ypredec1_xa_64x8m81_0/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_xa_64x8m81_6/a_n1_81# ypredec1_xa_64x8m81_5/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_xa_64x8m81_6/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_xa_64x8m81_7/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ a_6100_2150# ypredec1_xa_64x8m81_3/a_n1_81# a_975_1949# ypredec1_xa_64x8m81_4/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ a_6324_2352# ypredec1_xa_64x8m81_0/a_n1_81# ypredec1_xa_64x8m81_7/a_n1_81# ypredec1_xa_64x8m81_7/pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/S
+ ypredec1_xa_64x8m81_3/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ a_751_2554# a_303_2957# VSUBS
Xypredec1_xa_64x8m81_0 a_527_2758# a_6100_2150# a_975_1949# VSUBS a_6324_2352# a_751_2554#
+ a_303_2957# a_527_2758# ypredec1_xa_64x8m81_0/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_xa_64x8m81_0/a_n1_81# a_751_2554# a_6324_2352# ypredec1_xa_64x8m81_7/pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/S
+ VSUBS ypredec1_xa_64x8m81
Xypredec1_xa_64x8m81_1 a_527_2758# a_6100_2150# a_975_1949# VSUBS a_6324_2352# a_751_2554#
+ a_303_2957# a_6100_2150# ypredec1_xa_64x8m81_1/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ VSUBS a_751_2554# a_6324_2352# ypredec1_xa_64x8m81_7/pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/S
+ VSUBS ypredec1_xa_64x8m81
Xypredec1_xa_64x8m81_2 a_527_2758# a_6100_2150# a_975_1949# VSUBS a_303_2957# a_751_2554#
+ a_303_2957# a_6100_2150# ypredec1_xa_64x8m81_2/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ VSUBS a_751_2554# a_6324_2352# ypredec1_xa_64x8m81_7/pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/S
+ VSUBS ypredec1_xa_64x8m81
Xypredec1_xa_64x8m81_4 a_527_2758# a_6100_2150# a_975_1949# VSUBS a_6324_2352# a_751_2554#
+ a_303_2957# a_527_2758# ypredec1_xa_64x8m81_4/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_xa_64x8m81_4/a_n1_81# a_975_1949# a_6324_2352# ypredec1_xa_64x8m81_7/pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/S
+ VSUBS ypredec1_xa_64x8m81
Xypredec1_xa_64x8m81_3 a_527_2758# a_6100_2150# a_975_1949# VSUBS a_303_2957# a_751_2554#
+ a_303_2957# a_527_2758# ypredec1_xa_64x8m81_3/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_xa_64x8m81_3/a_n1_81# a_751_2554# a_6324_2352# ypredec1_xa_64x8m81_7/pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/S
+ VSUBS ypredec1_xa_64x8m81
Xypredec1_xa_64x8m81_5 a_527_2758# a_6100_2150# a_975_1949# VSUBS a_6324_2352# a_751_2554#
+ a_303_2957# a_6100_2150# ypredec1_xa_64x8m81_5/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ VSUBS a_975_1949# a_6324_2352# ypredec1_xa_64x8m81_7/pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/S
+ VSUBS ypredec1_xa_64x8m81
Xypredec1_xa_64x8m81_6 a_527_2758# a_6100_2150# a_975_1949# VSUBS a_303_2957# a_751_2554#
+ a_303_2957# a_6100_2150# ypredec1_xa_64x8m81_6/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_xa_64x8m81_6/a_n1_81# a_975_1949# a_6324_2352# ypredec1_xa_64x8m81_7/pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/S
+ VSUBS ypredec1_xa_64x8m81
Xypredec1_xa_64x8m81_7 a_527_2758# a_6100_2150# a_975_1949# VSUBS a_303_2957# a_751_2554#
+ a_303_2957# a_527_2758# ypredec1_xa_64x8m81_7/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_xa_64x8m81_7/a_n1_81# a_975_1949# a_6324_2352# ypredec1_xa_64x8m81_7/pmos_1p2$$47821868_64x8m81_2/pmos_5p04310589983264_64x8m81_0/S
+ VSUBS ypredec1_xa_64x8m81
.ends

.subckt pmos_5p04310589983259_64x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=20u l=0.6u
.ends

.subckt nmos_5p04310589983258_64x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=9.08u l=0.6u
.ends

.subckt ypredec1_ys_64x8m81 a_254_2184# nmos_5p04310589983258_64x8m81_1/D nmos_5p04310589983258_64x8m81_3/D
+ nmos_5p04310589983258_64x8m81_2/S pmos_5p04310589983259_64x8m81_3/S pmos_5p04310589983259_64x8m81_1/S
+ pmos_5p04310589983259_64x8m81_3/D VSUBS
Xpmos_5p04310589983259_64x8m81_2 pmos_5p04310589983259_64x8m81_3/D pmos_5p04310589983259_64x8m81_3/S
+ pmos_5p04310589983259_64x8m81_0/D pmos_5p04310589983259_64x8m81_3/D pmos_5p04310589983259_64x8m81
Xpmos_5p04310589983259_64x8m81_3 pmos_5p04310589983259_64x8m81_3/D pmos_5p04310589983259_64x8m81_3/D
+ pmos_5p04310589983259_64x8m81_0/D pmos_5p04310589983259_64x8m81_3/S pmos_5p04310589983259_64x8m81
Xnmos_5p04310589983258_64x8m81_0 pmos_5p04310589983259_64x8m81_3/S pmos_5p04310589983259_64x8m81_0/D
+ nmos_5p04310589983258_64x8m81_1/D VSUBS nmos_5p04310589983258_64x8m81
Xnmos_5p04310589983258_64x8m81_1 nmos_5p04310589983258_64x8m81_1/D pmos_5p04310589983259_64x8m81_0/D
+ pmos_5p04310589983259_64x8m81_1/S VSUBS nmos_5p04310589983258_64x8m81
Xnmos_5p04310589983258_64x8m81_2 pmos_5p04310589983259_64x8m81_0/D a_254_2184# nmos_5p04310589983258_64x8m81_2/S
+ VSUBS nmos_5p04310589983258_64x8m81
Xnmos_5p04310589983258_64x8m81_3 nmos_5p04310589983258_64x8m81_3/D pmos_5p04310589983259_64x8m81_0/D
+ pmos_5p04310589983259_64x8m81_3/S VSUBS nmos_5p04310589983258_64x8m81
Xpmos_5p04310589983259_64x8m81_0 pmos_5p04310589983259_64x8m81_3/D pmos_5p04310589983259_64x8m81_0/D
+ a_254_2184# pmos_5p04310589983259_64x8m81_3/D pmos_5p04310589983259_64x8m81
Xpmos_5p04310589983259_64x8m81_1 pmos_5p04310589983259_64x8m81_3/D pmos_5p04310589983259_64x8m81_3/D
+ pmos_5p04310589983259_64x8m81_0/D pmos_5p04310589983259_64x8m81_1/S pmos_5p04310589983259_64x8m81
.ends

.subckt pmos_5p04310589983266_64x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=1.71u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.71u l=0.6u
.ends

.subckt pmos_1p2$$47109164_64x8m81 a_n31_341# pmos_5p04310589983266_64x8m81_0/w_n208_n120#
+ pmos_5p04310589983266_64x8m81_0/S pmos_5p04310589983266_64x8m81_0/D a_193_341#
Xpmos_5p04310589983266_64x8m81_0 pmos_5p04310589983266_64x8m81_0/w_n208_n120# pmos_5p04310589983266_64x8m81_0/D
+ a_n31_341# pmos_5p04310589983266_64x8m81_0/S a_193_341# pmos_5p04310589983266_64x8m81
.ends

.subckt ypredec1_64x8m81 ly[5] ly[4] ly[7] ly[3] ly[2] ly[1] ly[0] ry[0] ry[1] ry[2]
+ ry[3] ry[4] ry[5] ry[6] ry[7] ly[6] men A[0] A[1] A[2] clk ypredec1_ys_64x8m81_9/pmos_5p04310589983259_64x8m81_3/D
+ ypredec1_bot_64x8m81_2/alatch_64x8m81_0/vdd ypredec1_ys_64x8m81_9/VSUBS pmos_1p2$$47109164_64x8m81_0/pmos_5p04310589983266_64x8m81_0/w_n208_n120#
+ ypredec1_bot_64x8m81_2/pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/S
+ pmos_1p2$$47109164_64x8m81_0/pmos_5p04310589983266_64x8m81_0/S
Xypredec1_bot_64x8m81_0 ypredec1_bot_64x8m81_2/pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/D
+ ypredec1_bot_64x8m81_2/pmos_1p2$$46887980_64x8m81_0/pmos_5p0431058998324_64x8m81_0/D
+ ypredec1_bot_64x8m81_2/pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/S
+ ypredec1_ys_64x8m81_9/VSUBS ypredec1_bot_64x8m81_1/pmos_1p2$$46887980_64x8m81_0/pmos_5p0431058998324_64x8m81_0/D
+ ypredec1_bot_64x8m81_2/alatch_64x8m81_0/enb ypredec1_bot_64x8m81_0/pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/D
+ ypredec1_bot_64x8m81_1/pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/D
+ ypredec1_bot_64x8m81_2/alatch_64x8m81_0/vdd ypredec1_bot_64x8m81_0/pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/D
+ ypredec1_bot_64x8m81_0/pmos_1p2$$46887980_64x8m81_0/pmos_5p0431058998324_64x8m81_0/D
+ A[0] ypredec1_bot_64x8m81_0/pmos_1p2$$46887980_64x8m81_0/pmos_5p0431058998324_64x8m81_0/D
+ nmos_5p04310589983260_64x8m81_1/D ypredec1_bot_64x8m81
Xypredec1_bot_64x8m81_1 ypredec1_bot_64x8m81_2/pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/D
+ ypredec1_bot_64x8m81_2/pmos_1p2$$46887980_64x8m81_0/pmos_5p0431058998324_64x8m81_0/D
+ ypredec1_bot_64x8m81_2/pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/S
+ ypredec1_ys_64x8m81_9/VSUBS ypredec1_bot_64x8m81_1/pmos_1p2$$46887980_64x8m81_0/pmos_5p0431058998324_64x8m81_0/D
+ ypredec1_bot_64x8m81_2/alatch_64x8m81_0/enb ypredec1_bot_64x8m81_0/pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/D
+ ypredec1_bot_64x8m81_1/pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/D
+ ypredec1_bot_64x8m81_2/alatch_64x8m81_0/vdd ypredec1_bot_64x8m81_1/pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/D
+ ypredec1_bot_64x8m81_0/pmos_1p2$$46887980_64x8m81_0/pmos_5p0431058998324_64x8m81_0/D
+ A[2] ypredec1_bot_64x8m81_1/pmos_1p2$$46887980_64x8m81_0/pmos_5p0431058998324_64x8m81_0/D
+ nmos_5p04310589983260_64x8m81_1/D ypredec1_bot_64x8m81
Xypredec1_bot_64x8m81_2 ypredec1_bot_64x8m81_2/pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/D
+ ypredec1_bot_64x8m81_2/pmos_1p2$$46887980_64x8m81_0/pmos_5p0431058998324_64x8m81_0/D
+ ypredec1_bot_64x8m81_2/pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/S
+ ypredec1_ys_64x8m81_9/VSUBS ypredec1_bot_64x8m81_1/pmos_1p2$$46887980_64x8m81_0/pmos_5p0431058998324_64x8m81_0/D
+ ypredec1_bot_64x8m81_2/alatch_64x8m81_0/enb ypredec1_bot_64x8m81_0/pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/D
+ ypredec1_bot_64x8m81_1/pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/D
+ ypredec1_bot_64x8m81_2/alatch_64x8m81_0/vdd ypredec1_bot_64x8m81_2/pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/D
+ ypredec1_bot_64x8m81_0/pmos_1p2$$46887980_64x8m81_0/pmos_5p0431058998324_64x8m81_0/D
+ A[1] ypredec1_bot_64x8m81_2/pmos_1p2$$46887980_64x8m81_0/pmos_5p0431058998324_64x8m81_0/D
+ nmos_5p04310589983260_64x8m81_1/D ypredec1_bot_64x8m81
Xnmos_5p04310589983260_64x8m81_0 ypredec1_ys_64x8m81_9/VSUBS clk nmos_5p04310589983260_64x8m81_1/D
+ ypredec1_ys_64x8m81_9/VSUBS nmos_5p04310589983260_64x8m81
Xnmos_5p04310589983260_64x8m81_1 nmos_5p04310589983260_64x8m81_1/D men ypredec1_ys_64x8m81_9/VSUBS
+ ypredec1_ys_64x8m81_9/VSUBS nmos_5p04310589983260_64x8m81
Xypredec1_xax8_64x8m81_0 ypredec1_xax8_64x8m81_0/ypredec1_xa_64x8m81_1/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_xax8_64x8m81_0/ypredec1_xa_64x8m81_2/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_bot_64x8m81_2/pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/D
+ ypredec1_xax8_64x8m81_0/ypredec1_xa_64x8m81_0/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_ys_64x8m81_9/VSUBS ypredec1_xax8_64x8m81_0/ypredec1_xa_64x8m81_5/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_xax8_64x8m81_0/ypredec1_xa_64x8m81_6/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_xax8_64x8m81_0/ypredec1_xa_64x8m81_7/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_bot_64x8m81_2/pmos_1p2$$46887980_64x8m81_0/pmos_5p0431058998324_64x8m81_0/D
+ ypredec1_ys_64x8m81_9/VSUBS ypredec1_bot_64x8m81_0/pmos_1p2$$46887980_64x8m81_0/pmos_5p0431058998324_64x8m81_0/D
+ ypredec1_xax8_64x8m81_0/ypredec1_xa_64x8m81_4/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_bot_64x8m81_1/pmos_1p2$$46887980_64x8m81_0/pmos_5p0431058998324_64x8m81_0/D
+ ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS ypredec1_bot_64x8m81_2/pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/S
+ ypredec1_xax8_64x8m81_0/ypredec1_xa_64x8m81_3/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_bot_64x8m81_0/pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/D
+ ypredec1_bot_64x8m81_1/pmos_1p2$$46887980_64x8m81_1/pmos_5p0431058998324_64x8m81_0/D
+ ypredec1_ys_64x8m81_9/VSUBS ypredec1_xax8_64x8m81
Xypredec1_ys_64x8m81_10 ypredec1_xax8_64x8m81_0/ypredec1_xa_64x8m81_6/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS
+ ry[4] ry[4] ypredec1_ys_64x8m81_9/pmos_5p04310589983259_64x8m81_3/D ypredec1_ys_64x8m81_9/VSUBS
+ ypredec1_ys_64x8m81
Xypredec1_ys_64x8m81_11 ypredec1_xax8_64x8m81_0/ypredec1_xa_64x8m81_2/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS
+ ry[5] ry[5] ypredec1_ys_64x8m81_9/pmos_5p04310589983259_64x8m81_3/D ypredec1_ys_64x8m81_9/VSUBS
+ ypredec1_ys_64x8m81
Xypredec1_ys_64x8m81_12 ypredec1_xax8_64x8m81_0/ypredec1_xa_64x8m81_7/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS
+ ry[6] ry[6] ypredec1_ys_64x8m81_9/pmos_5p04310589983259_64x8m81_3/D ypredec1_ys_64x8m81_9/VSUBS
+ ypredec1_ys_64x8m81
Xypredec1_ys_64x8m81_13 ypredec1_xax8_64x8m81_0/ypredec1_xa_64x8m81_3/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS
+ ry[7] ry[7] ypredec1_ys_64x8m81_9/pmos_5p04310589983259_64x8m81_3/D ypredec1_ys_64x8m81_9/VSUBS
+ ypredec1_ys_64x8m81
Xypredec1_ys_64x8m81_14 ypredec1_xax8_64x8m81_0/ypredec1_xa_64x8m81_5/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS
+ ry[0] ry[0] ypredec1_ys_64x8m81_9/pmos_5p04310589983259_64x8m81_3/D ypredec1_ys_64x8m81_9/VSUBS
+ ypredec1_ys_64x8m81
Xypredec1_ys_64x8m81_15 ypredec1_xax8_64x8m81_0/ypredec1_xa_64x8m81_3/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS
+ ly[7] ly[7] ypredec1_ys_64x8m81_9/pmos_5p04310589983259_64x8m81_3/D ypredec1_ys_64x8m81_9/VSUBS
+ ypredec1_ys_64x8m81
Xnmos_1p2$$47342636_64x8m81_0 ypredec1_bot_64x8m81_2/alatch_64x8m81_0/enb ypredec1_ys_64x8m81_9/VSUBS
+ nmos_5p04310589983260_64x8m81_1/D ypredec1_ys_64x8m81_9/VSUBS nmos_1p2$$47342636_64x8m81
Xypredec1_ys_64x8m81_0 ypredec1_xax8_64x8m81_0/ypredec1_xa_64x8m81_5/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS
+ ly[0] ly[0] ypredec1_ys_64x8m81_9/pmos_5p04310589983259_64x8m81_3/D ypredec1_ys_64x8m81_9/VSUBS
+ ypredec1_ys_64x8m81
Xypredec1_ys_64x8m81_1 ypredec1_xax8_64x8m81_0/ypredec1_xa_64x8m81_1/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS
+ ly[1] ly[1] ypredec1_ys_64x8m81_9/pmos_5p04310589983259_64x8m81_3/D ypredec1_ys_64x8m81_9/VSUBS
+ ypredec1_ys_64x8m81
Xypredec1_ys_64x8m81_2 ypredec1_xax8_64x8m81_0/ypredec1_xa_64x8m81_4/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS
+ ly[2] ly[2] ypredec1_ys_64x8m81_9/pmos_5p04310589983259_64x8m81_3/D ypredec1_ys_64x8m81_9/VSUBS
+ ypredec1_ys_64x8m81
Xypredec1_ys_64x8m81_3 ypredec1_xax8_64x8m81_0/ypredec1_xa_64x8m81_0/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS
+ ly[3] ly[3] ypredec1_ys_64x8m81_9/pmos_5p04310589983259_64x8m81_3/D ypredec1_ys_64x8m81_9/VSUBS
+ ypredec1_ys_64x8m81
Xypredec1_ys_64x8m81_4 ypredec1_xax8_64x8m81_0/ypredec1_xa_64x8m81_6/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS
+ ly[4] ly[4] ypredec1_ys_64x8m81_9/pmos_5p04310589983259_64x8m81_3/D ypredec1_ys_64x8m81_9/VSUBS
+ ypredec1_ys_64x8m81
Xypredec1_ys_64x8m81_5 ypredec1_xax8_64x8m81_0/ypredec1_xa_64x8m81_2/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS
+ ly[5] ly[5] ypredec1_ys_64x8m81_9/pmos_5p04310589983259_64x8m81_3/D ypredec1_ys_64x8m81_9/VSUBS
+ ypredec1_ys_64x8m81
Xypredec1_ys_64x8m81_6 ypredec1_xax8_64x8m81_0/ypredec1_xa_64x8m81_7/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS
+ ly[6] ly[6] ypredec1_ys_64x8m81_9/pmos_5p04310589983259_64x8m81_3/D ypredec1_ys_64x8m81_9/VSUBS
+ ypredec1_ys_64x8m81
Xypredec1_ys_64x8m81_7 ypredec1_xax8_64x8m81_0/ypredec1_xa_64x8m81_1/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS
+ ry[1] ry[1] ypredec1_ys_64x8m81_9/pmos_5p04310589983259_64x8m81_3/D ypredec1_ys_64x8m81_9/VSUBS
+ ypredec1_ys_64x8m81
Xypredec1_ys_64x8m81_8 ypredec1_xax8_64x8m81_0/ypredec1_xa_64x8m81_4/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS
+ ry[2] ry[2] ypredec1_ys_64x8m81_9/pmos_5p04310589983259_64x8m81_3/D ypredec1_ys_64x8m81_9/VSUBS
+ ypredec1_ys_64x8m81
Xypredec1_ys_64x8m81_9 ypredec1_xax8_64x8m81_0/ypredec1_xa_64x8m81_0/nmos_1p2$$46551084_64x8m81_2/nmos_5p0431058998325_64x8m81_0/D
+ ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS ypredec1_ys_64x8m81_9/VSUBS
+ ry[3] ry[3] ypredec1_ys_64x8m81_9/pmos_5p04310589983259_64x8m81_3/D ypredec1_ys_64x8m81_9/VSUBS
+ ypredec1_ys_64x8m81
Xpmos_1p2$$47109164_64x8m81_0 nmos_5p04310589983260_64x8m81_1/D pmos_1p2$$47109164_64x8m81_0/pmos_5p04310589983266_64x8m81_0/w_n208_n120#
+ pmos_1p2$$47109164_64x8m81_0/pmos_5p04310589983266_64x8m81_0/S ypredec1_bot_64x8m81_2/alatch_64x8m81_0/enb
+ nmos_5p04310589983260_64x8m81_1/D pmos_1p2$$47109164_64x8m81
X0 a_7843_267# clk nmos_5p04310589983260_64x8m81_1/D pmos_1p2$$47109164_64x8m81_0/pmos_5p04310589983266_64x8m81_0/S pmos_3p3 w=2.275u l=0.6u
X1 nmos_5p04310589983260_64x8m81_1/D clk a_7395_267# pmos_1p2$$47109164_64x8m81_0/pmos_5p04310589983266_64x8m81_0/S pmos_3p3 w=2.275u l=0.6u
X2 a_7395_267# men pmos_1p2$$47109164_64x8m81_0/pmos_5p04310589983266_64x8m81_0/S pmos_1p2$$47109164_64x8m81_0/pmos_5p04310589983266_64x8m81_0/S pmos_3p3 w=2.275u l=0.6u
X3 pmos_1p2$$47109164_64x8m81_0/pmos_5p04310589983266_64x8m81_0/S men a_7843_267# pmos_1p2$$47109164_64x8m81_0/pmos_5p04310589983266_64x8m81_0/S pmos_3p3 w=2.275u l=0.6u
.ends

.subckt pmos_5p04310589983276_64x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=10.43u l=0.6u
.ends

.subckt pmos_1p2$$47512620_64x8m81 pmos_5p04310589983276_64x8m81_0/S a_n30_n74# pmos_5p04310589983276_64x8m81_0/D
+ w_n286_n142#
Xpmos_5p04310589983276_64x8m81_0 w_n286_n142# pmos_5p04310589983276_64x8m81_0/D a_n30_n74#
+ pmos_5p04310589983276_64x8m81_0/S pmos_5p04310589983276_64x8m81
.ends

.subckt pmos_5p04310589983272_64x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=11.34u l=0.6u
.ends

.subckt pmos_1p2$$47513644_64x8m81 pmos_5p04310589983272_64x8m81_0/S a_n30_n74# pmos_5p04310589983272_64x8m81_0/D
+ w_n286_n141#
Xpmos_5p04310589983272_64x8m81_0 w_n286_n141# pmos_5p04310589983272_64x8m81_0/D a_n30_n74#
+ pmos_5p04310589983272_64x8m81_0/S pmos_5p04310589983272_64x8m81
.ends

.subckt xpredec1_xa_64x8m81 a_197_n10255# m1_n58_n7539# a_421_n10255# m1_n58_n6933#
+ a_645_n10255# m1_n58_n7135# m1_n58_n6530# m1_n58_n7337# a_n1_81# pmos_1p2$$47513644_64x8m81_2/pmos_5p04310589983272_64x8m81_0/D
+ m1_n58_n6732# pmos_1p2$$47513644_64x8m81_2/pmos_5p04310589983272_64x8m81_0/S M3_M2$$47333420_64x8m81_1/VSUBS
Xpmos_1p2$$47512620_64x8m81_0 pmos_1p2$$47513644_64x8m81_2/pmos_5p04310589983272_64x8m81_0/S
+ a_645_n10255# pmos_1p2$$47512620_64x8m81_2/pmos_5p04310589983276_64x8m81_0/D pmos_1p2$$47513644_64x8m81_2/pmos_5p04310589983272_64x8m81_0/S
+ pmos_1p2$$47512620_64x8m81
Xpmos_1p2$$47513644_64x8m81_0 pmos_1p2$$47513644_64x8m81_2/pmos_5p04310589983272_64x8m81_0/D
+ pmos_1p2$$47512620_64x8m81_2/pmos_5p04310589983276_64x8m81_0/D pmos_1p2$$47513644_64x8m81_2/pmos_5p04310589983272_64x8m81_0/S
+ pmos_1p2$$47513644_64x8m81_2/pmos_5p04310589983272_64x8m81_0/S pmos_1p2$$47513644_64x8m81
Xpmos_1p2$$47512620_64x8m81_2 pmos_1p2$$47513644_64x8m81_2/pmos_5p04310589983272_64x8m81_0/S
+ a_197_n10255# pmos_1p2$$47512620_64x8m81_2/pmos_5p04310589983276_64x8m81_0/D pmos_1p2$$47513644_64x8m81_2/pmos_5p04310589983272_64x8m81_0/S
+ pmos_1p2$$47512620_64x8m81
Xpmos_1p2$$47512620_64x8m81_1 pmos_1p2$$47512620_64x8m81_2/pmos_5p04310589983276_64x8m81_0/D
+ a_421_n10255# pmos_1p2$$47513644_64x8m81_2/pmos_5p04310589983272_64x8m81_0/S pmos_1p2$$47513644_64x8m81_2/pmos_5p04310589983272_64x8m81_0/S
+ pmos_1p2$$47512620_64x8m81
Xpmos_1p2$$47513644_64x8m81_1 pmos_1p2$$47513644_64x8m81_2/pmos_5p04310589983272_64x8m81_0/S
+ pmos_1p2$$47512620_64x8m81_2/pmos_5p04310589983276_64x8m81_0/D pmos_1p2$$47513644_64x8m81_2/pmos_5p04310589983272_64x8m81_0/D
+ pmos_1p2$$47513644_64x8m81_2/pmos_5p04310589983272_64x8m81_0/S pmos_1p2$$47513644_64x8m81
Xpmos_1p2$$47513644_64x8m81_2 pmos_1p2$$47513644_64x8m81_2/pmos_5p04310589983272_64x8m81_0/S
+ pmos_1p2$$47512620_64x8m81_2/pmos_5p04310589983276_64x8m81_0/D pmos_1p2$$47513644_64x8m81_2/pmos_5p04310589983272_64x8m81_0/D
+ pmos_1p2$$47513644_64x8m81_2/pmos_5p04310589983272_64x8m81_0/S pmos_1p2$$47513644_64x8m81
Xnmos_1p2$$47514668_64x8m81_0 pmos_1p2$$47513644_64x8m81_2/pmos_5p04310589983272_64x8m81_0/D
+ pmos_1p2$$47512620_64x8m81_2/pmos_5p04310589983276_64x8m81_0/D M3_M2$$47333420_64x8m81_1/VSUBS
+ M3_M2$$47333420_64x8m81_1/VSUBS nmos_1p2$$47514668_64x8m81
Xnmos_1p2$$47514668_64x8m81_1 M3_M2$$47333420_64x8m81_1/VSUBS pmos_1p2$$47512620_64x8m81_2/pmos_5p04310589983276_64x8m81_0/D
+ pmos_1p2$$47513644_64x8m81_2/pmos_5p04310589983272_64x8m81_0/D M3_M2$$47333420_64x8m81_1/VSUBS
+ nmos_1p2$$47514668_64x8m81
Xnmos_1p2$$47514668_64x8m81_2 pmos_1p2$$47513644_64x8m81_2/pmos_5p04310589983272_64x8m81_0/D
+ pmos_1p2$$47512620_64x8m81_2/pmos_5p04310589983276_64x8m81_0/D M3_M2$$47333420_64x8m81_1/VSUBS
+ M3_M2$$47333420_64x8m81_1/VSUBS nmos_1p2$$47514668_64x8m81
X0 pmos_1p2$$47512620_64x8m81_2/pmos_5p04310589983276_64x8m81_0/D a_645_n10255# a_541_n10182# M3_M2$$47333420_64x8m81_1/VSUBS nmos_3p3 w=12.475u l=0.6u
X1 a_317_n10182# a_197_n10255# M3_M2$$47333420_64x8m81_1/VSUBS M3_M2$$47333420_64x8m81_1/VSUBS nmos_3p3 w=12.475u l=0.6u
X2 a_541_n10182# a_421_n10255# a_317_n10182# M3_M2$$47333420_64x8m81_1/VSUBS nmos_3p3 w=12.475u l=0.6u
.ends

.subckt nmos_5p04310589983275_64x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=6.58u l=0.6u
.ends

.subckt nmos_1p2$$47336492_64x8m81 nmos_5p04310589983275_64x8m81_0/D nmos_5p04310589983275_64x8m81_0/S
+ a_n31_n74# VSUBS
Xnmos_5p04310589983275_64x8m81_0 nmos_5p04310589983275_64x8m81_0/D a_n31_n74# nmos_5p04310589983275_64x8m81_0/S
+ VSUBS nmos_5p04310589983275_64x8m81
.ends

.subckt pmos_5p04310589983274_64x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=16.33u l=0.6u
.ends

.subckt pmos_1p2$$47337516_64x8m81 pmos_5p04310589983274_64x8m81_0/S pmos_5p04310589983274_64x8m81_0/D
+ a_n31_n73# w_n286_n141#
Xpmos_5p04310589983274_64x8m81_0 w_n286_n141# pmos_5p04310589983274_64x8m81_0/D a_n31_n73#
+ pmos_5p04310589983274_64x8m81_0/S pmos_5p04310589983274_64x8m81
.ends

.subckt xpredec1_bot_64x8m81 m1_n106_2472# m1_n106_3279# m1_n106_2674# alatch_64x8m81_0/enb
+ alatch_64x8m81_0/vdd pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/S m1_n106_2876# alatch_64x8m81_0/a
+ pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D m1_n106_3078# m1_n106_3481#
+ VSUBS alatch_64x8m81_0/en
Xnmos_1p2$$47336492_64x8m81_0 pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ VSUBS pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D VSUBS nmos_1p2$$47336492_64x8m81
Xnmos_1p2$$47336492_64x8m81_1 pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ VSUBS alatch_64x8m81_0/ab VSUBS nmos_1p2$$47336492_64x8m81
Xalatch_64x8m81_0 alatch_64x8m81_0/enb alatch_64x8m81_0/en alatch_64x8m81_0/ab alatch_64x8m81_0/a
+ VSUBS alatch_64x8m81_0/vdd alatch_64x8m81
Xpmos_1p2$$47337516_64x8m81_0 pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/S
+ pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/S pmos_1p2$$47337516_64x8m81
Xpmos_1p2$$47337516_64x8m81_1 pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/S
+ pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D alatch_64x8m81_0/ab
+ pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/S pmos_1p2$$47337516_64x8m81
.ends

.subckt xpredec1_64x8m81 A[2] men x[7] x[6] x[5] x[4] x[3] x[2] x[1] x[0] A[1] A[0]
+ clk w_7178_9364# vdd pmos_1p2$$47109164_64x8m81_0/pmos_5p04310589983266_64x8m81_0/w_n208_n120#
+ vss
Xxpredec1_xa_64x8m81_4 xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ vss x[2] xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ vdd vss xpredec1_xa_64x8m81
Xxpredec1_xa_64x8m81_5 xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ vss x[0] xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ vdd vss xpredec1_xa_64x8m81
Xxpredec1_xa_64x8m81_6 xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ vss x[4] xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ vdd vss xpredec1_xa_64x8m81
Xxpredec1_xa_64x8m81_7 xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_xa_64x8m81_7/a_n1_81# x[6] xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ vdd vss xpredec1_xa_64x8m81
Xnmos_5p04310589983260_64x8m81_0 vss clk nmos_5p04310589983260_64x8m81_1/D vss nmos_5p04310589983260_64x8m81
Xnmos_5p04310589983260_64x8m81_1 nmos_5p04310589983260_64x8m81_1/D men vss vss nmos_5p04310589983260_64x8m81
Xnmos_1p2$$47342636_64x8m81_0 xpredec1_bot_64x8m81_2/alatch_64x8m81_0/enb vss nmos_5p04310589983260_64x8m81_1/D
+ vss nmos_1p2$$47342636_64x8m81
Xxpredec1_bot_64x8m81_0 xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_2/alatch_64x8m81_0/enb vdd xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ vdd xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ A[0] xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ vss nmos_5p04310589983260_64x8m81_1/D xpredec1_bot_64x8m81
Xxpredec1_bot_64x8m81_1 xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_2/alatch_64x8m81_0/enb vdd xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ vdd xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ A[2] xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ vss nmos_5p04310589983260_64x8m81_1/D xpredec1_bot_64x8m81
Xxpredec1_bot_64x8m81_2 xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_2/alatch_64x8m81_0/enb vdd xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ vdd xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ A[1] xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ vss nmos_5p04310589983260_64x8m81_1/D xpredec1_bot_64x8m81
Xxpredec1_xa_64x8m81_0 xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ vss x[3] xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ vdd vss xpredec1_xa_64x8m81
Xxpredec1_xa_64x8m81_1 xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_xa_64x8m81_1/a_n1_81# x[1] xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ vdd vss xpredec1_xa_64x8m81
Xpmos_1p2$$47109164_64x8m81_0 nmos_5p04310589983260_64x8m81_1/D pmos_1p2$$47109164_64x8m81_0/pmos_5p04310589983266_64x8m81_0/w_n208_n120#
+ vdd xpredec1_bot_64x8m81_2/alatch_64x8m81_0/enb nmos_5p04310589983260_64x8m81_1/D
+ pmos_1p2$$47109164_64x8m81
Xxpredec1_xa_64x8m81_2 xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ vss x[5] xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ vdd vss xpredec1_xa_64x8m81
Xxpredec1_xa_64x8m81_3 xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_0/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_1/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_0/pmos_5p04310589983274_64x8m81_0/D
+ xpredec1_xa_64x8m81_3/a_n1_81# x[7] xpredec1_bot_64x8m81_2/pmos_1p2$$47337516_64x8m81_1/pmos_5p04310589983274_64x8m81_0/D
+ vdd vss xpredec1_xa_64x8m81
X0 nmos_5p04310589983260_64x8m81_1/D clk a_7553_9505# w_7178_9364# pmos_3p3 w=2.275u l=0.6u
X1 a_7553_9505# men vdd w_7178_9364# pmos_3p3 w=2.275u l=0.6u
X2 a_8001_9505# clk nmos_5p04310589983260_64x8m81_1/D w_7178_9364# pmos_3p3 w=2.275u l=0.6u
X3 vdd men a_8001_9505# w_7178_9364# pmos_3p3 w=2.275u l=0.6u
.ends

.subckt pmos_5p04310589983268_64x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=17.69u l=0.6u
.ends

.subckt pmos_1p2$$47503404_64x8m81 a_n31_n73# pmos_5p04310589983268_64x8m81_0/S w_n286_n141#
+ pmos_5p04310589983268_64x8m81_0/D
Xpmos_5p04310589983268_64x8m81_0 w_n286_n141# pmos_5p04310589983268_64x8m81_0/D a_n31_n73#
+ pmos_5p04310589983268_64x8m81_0/S pmos_5p04310589983268_64x8m81
.ends

.subckt nmos_5p04310589983270_64x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=7.04u l=0.6u
.ends

.subckt pmos_5p04310589983267_64x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=13.16u l=0.6u
.ends

.subckt pmos_1p2$$47504428_64x8m81 pmos_5p04310589983267_64x8m81_0/S w_n286_n142#
+ pmos_5p04310589983267_64x8m81_0/w_n208_n120# a_n31_n73# pmos_5p04310589983267_64x8m81_0/D
Xpmos_5p04310589983267_64x8m81_0 pmos_5p04310589983267_64x8m81_0/w_n208_n120# pmos_5p04310589983267_64x8m81_0/D
+ a_n31_n73# pmos_5p04310589983267_64x8m81_0/S pmos_5p04310589983267_64x8m81
.ends

.subckt nmos_5p04310589983269_64x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=5.22u l=0.6u
.ends

.subckt nmos_1p2$$47502380_64x8m81 nmos_5p04310589983269_64x8m81_0/D a_n31_n74# VSUBS
+ nmos_5p04310589983269_64x8m81_0/S
Xnmos_5p04310589983269_64x8m81_0 nmos_5p04310589983269_64x8m81_0/D a_n31_n74# nmos_5p04310589983269_64x8m81_0/S
+ VSUBS nmos_5p04310589983269_64x8m81
.ends

.subckt xpredec0_bot_64x8m81 m1_n106_2472# m1_n106_2674# alatch_64x8m81_0/enb alatch_64x8m81_0/vdd
+ pmos_1p2$$47504428_64x8m81_0/pmos_5p04310589983267_64x8m81_0/D nmos_5p04310589983270_64x8m81_0/D
+ m1_n106_2876# alatch_64x8m81_0/a pmos_1p2$$47504428_64x8m81_0/pmos_5p04310589983267_64x8m81_0/S
+ m1_n106_3078# VSUBS alatch_64x8m81_0/en
Xpmos_1p2$$47503404_64x8m81_0 alatch_64x8m81_0/ab pmos_1p2$$47504428_64x8m81_0/pmos_5p04310589983267_64x8m81_0/S
+ pmos_1p2$$47504428_64x8m81_0/pmos_5p04310589983267_64x8m81_0/S nmos_5p04310589983270_64x8m81_0/D
+ pmos_1p2$$47503404_64x8m81
Xnmos_5p04310589983270_64x8m81_0 nmos_5p04310589983270_64x8m81_0/D alatch_64x8m81_0/ab
+ VSUBS VSUBS nmos_5p04310589983270_64x8m81
Xpmos_1p2$$47504428_64x8m81_0 pmos_1p2$$47504428_64x8m81_0/pmos_5p04310589983267_64x8m81_0/S
+ pmos_1p2$$47504428_64x8m81_0/pmos_5p04310589983267_64x8m81_0/S pmos_1p2$$47504428_64x8m81_0/pmos_5p04310589983267_64x8m81_0/S
+ nmos_5p04310589983270_64x8m81_0/D pmos_1p2$$47504428_64x8m81_0/pmos_5p04310589983267_64x8m81_0/D
+ pmos_1p2$$47504428_64x8m81
Xalatch_64x8m81_0 alatch_64x8m81_0/enb alatch_64x8m81_0/en alatch_64x8m81_0/ab alatch_64x8m81_0/a
+ VSUBS alatch_64x8m81_0/vdd alatch_64x8m81
Xnmos_1p2$$47502380_64x8m81_0 pmos_1p2$$47504428_64x8m81_0/pmos_5p04310589983267_64x8m81_0/D
+ nmos_5p04310589983270_64x8m81_0/D VSUBS VSUBS nmos_1p2$$47502380_64x8m81
.ends

.subckt pmos_5p04310589983273_64x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=1.14u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.14u l=0.6u
.ends

.subckt nmos_5p04310589983240_64x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=1.37u l=0.6u
.ends

.subckt pmos_5p04310589983271_64x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=15.2u l=0.6u
.ends

.subckt pmos_1p2$$47643692_64x8m81 pmos_5p04310589983271_64x8m81_0/S pmos_5p04310589983271_64x8m81_0/D
+ w_n286_n142# a_n31_n74#
Xpmos_5p04310589983271_64x8m81_0 w_n286_n142# pmos_5p04310589983271_64x8m81_0/D a_n31_n74#
+ pmos_5p04310589983271_64x8m81_0/S pmos_5p04310589983271_64x8m81
.ends

.subckt nmos_1p2$$47641644_64x8m81 a_n31_n73# nmos_5p04310589983261_64x8m81_0/D nmos_5p04310589983261_64x8m81_0/S
+ VSUBS
Xnmos_5p04310589983261_64x8m81_0 nmos_5p04310589983261_64x8m81_0/D a_n31_n73# nmos_5p04310589983261_64x8m81_0/S
+ VSUBS nmos_5p04310589983261_64x8m81
.ends

.subckt pmos_1p2$$47642668_64x8m81 pmos_5p04310589983271_64x8m81_0/S w_n546_n142#
+ pmos_5p04310589983271_64x8m81_0/D a_n31_n74#
Xpmos_5p04310589983271_64x8m81_0 w_n546_n142# pmos_5p04310589983271_64x8m81_0/D a_n31_n74#
+ pmos_5p04310589983271_64x8m81_0/S pmos_5p04310589983271_64x8m81
.ends

.subckt xpredec0_xa_64x8m81 nmos_1p2$$47641644_64x8m81_0/nmos_5p04310589983261_64x8m81_0/S
+ m1_342_3273# a_875_414# m3_855_1044# a_651_414# m1_342_3474# m3_153_8117# pmos_1p2$$47513644_64x8m81_3/pmos_5p04310589983272_64x8m81_0/D
+ m1_342_3071# m1_342_3676# pmos_1p2$$47513644_64x8m81_3/pmos_5p04310589983272_64x8m81_0/S
+ nmos_1p2$$47641644_64x8m81_3/nmos_5p04310589983261_64x8m81_0/D M3_M2$$47644716_64x8m81_2/VSUBS
+ pmos_1p2$$47643692_64x8m81_0/pmos_5p04310589983271_64x8m81_0/D
Xpmos_1p2$$47643692_64x8m81_0 pmos_1p2$$47643692_64x8m81_0/pmos_5p04310589983271_64x8m81_0/S
+ pmos_1p2$$47643692_64x8m81_0/pmos_5p04310589983271_64x8m81_0/D pmos_1p2$$47643692_64x8m81_0/pmos_5p04310589983271_64x8m81_0/D
+ a_651_414# pmos_1p2$$47643692_64x8m81
Xnmos_1p2$$47641644_64x8m81_2 pmos_1p2$$47643692_64x8m81_0/pmos_5p04310589983271_64x8m81_0/S
+ nmos_1p2$$47641644_64x8m81_3/nmos_5p04310589983261_64x8m81_0/D pmos_1p2$$47513644_64x8m81_3/pmos_5p04310589983272_64x8m81_0/D
+ M3_M2$$47644716_64x8m81_2/VSUBS nmos_1p2$$47641644_64x8m81
Xnmos_1p2$$47641644_64x8m81_3 pmos_1p2$$47643692_64x8m81_0/pmos_5p04310589983271_64x8m81_0/S
+ nmos_1p2$$47641644_64x8m81_3/nmos_5p04310589983261_64x8m81_0/D pmos_1p2$$47513644_64x8m81_3/pmos_5p04310589983272_64x8m81_0/D
+ M3_M2$$47644716_64x8m81_2/VSUBS nmos_1p2$$47641644_64x8m81
Xpmos_1p2$$47513644_64x8m81_0 pmos_1p2$$47513644_64x8m81_3/pmos_5p04310589983272_64x8m81_0/D
+ pmos_1p2$$47643692_64x8m81_0/pmos_5p04310589983271_64x8m81_0/S pmos_1p2$$47513644_64x8m81_3/pmos_5p04310589983272_64x8m81_0/S
+ pmos_1p2$$47643692_64x8m81_0/pmos_5p04310589983271_64x8m81_0/D pmos_1p2$$47513644_64x8m81
Xpmos_1p2$$47513644_64x8m81_1 pmos_1p2$$47513644_64x8m81_3/pmos_5p04310589983272_64x8m81_0/S
+ pmos_1p2$$47643692_64x8m81_0/pmos_5p04310589983271_64x8m81_0/S pmos_1p2$$47513644_64x8m81_3/pmos_5p04310589983272_64x8m81_0/D
+ pmos_1p2$$47643692_64x8m81_0/pmos_5p04310589983271_64x8m81_0/D pmos_1p2$$47513644_64x8m81
Xpmos_1p2$$47513644_64x8m81_2 pmos_1p2$$47513644_64x8m81_3/pmos_5p04310589983272_64x8m81_0/D
+ pmos_1p2$$47643692_64x8m81_0/pmos_5p04310589983271_64x8m81_0/S pmos_1p2$$47513644_64x8m81_3/pmos_5p04310589983272_64x8m81_0/S
+ pmos_1p2$$47643692_64x8m81_0/pmos_5p04310589983271_64x8m81_0/D pmos_1p2$$47513644_64x8m81
Xpmos_1p2$$47513644_64x8m81_3 pmos_1p2$$47513644_64x8m81_3/pmos_5p04310589983272_64x8m81_0/S
+ pmos_1p2$$47643692_64x8m81_0/pmos_5p04310589983271_64x8m81_0/S pmos_1p2$$47513644_64x8m81_3/pmos_5p04310589983272_64x8m81_0/D
+ pmos_1p2$$47643692_64x8m81_0/pmos_5p04310589983271_64x8m81_0/D pmos_1p2$$47513644_64x8m81
Xpmos_1p2$$47642668_64x8m81_0 pmos_1p2$$47643692_64x8m81_0/pmos_5p04310589983271_64x8m81_0/D
+ pmos_1p2$$47643692_64x8m81_0/pmos_5p04310589983271_64x8m81_0/D pmos_1p2$$47643692_64x8m81_0/pmos_5p04310589983271_64x8m81_0/S
+ a_875_414# pmos_1p2$$47642668_64x8m81
Xnmos_1p2$$47641644_64x8m81_0 pmos_1p2$$47643692_64x8m81_0/pmos_5p04310589983271_64x8m81_0/S
+ pmos_1p2$$47513644_64x8m81_3/pmos_5p04310589983272_64x8m81_0/D nmos_1p2$$47641644_64x8m81_0/nmos_5p04310589983261_64x8m81_0/S
+ M3_M2$$47644716_64x8m81_2/VSUBS nmos_1p2$$47641644_64x8m81
Xnmos_1p2$$47641644_64x8m81_1 pmos_1p2$$47643692_64x8m81_0/pmos_5p04310589983271_64x8m81_0/S
+ pmos_1p2$$47513644_64x8m81_3/pmos_5p04310589983272_64x8m81_0/D nmos_1p2$$47641644_64x8m81_3/nmos_5p04310589983261_64x8m81_0/D
+ M3_M2$$47644716_64x8m81_2/VSUBS nmos_1p2$$47641644_64x8m81
X0 a_771_486# a_651_414# pmos_1p2$$47643692_64x8m81_0/pmos_5p04310589983271_64x8m81_0/S M3_M2$$47644716_64x8m81_2/VSUBS nmos_3p3 w=12.25u l=0.6u
X1 M3_M2$$47644716_64x8m81_2/VSUBS a_875_414# a_771_486# M3_M2$$47644716_64x8m81_2/VSUBS nmos_3p3 w=12.25u l=0.6u
.ends

.subckt xpredec0_64x8m81 A[0] men x[0] x[1] x[2] x[3] A[1] clk xpredec0_xa_64x8m81_2/nmos_1p2$$47641644_64x8m81_0/nmos_5p04310589983261_64x8m81_0/S
+ xpredec0_xa_64x8m81_3/nmos_1p2$$47641644_64x8m81_0/nmos_5p04310589983261_64x8m81_0/S
+ vss vdd
Xxpredec0_bot_64x8m81_0 xpredec0_bot_64x8m81_0/pmos_1p2$$47504428_64x8m81_0/pmos_5p04310589983267_64x8m81_0/D
+ xpredec0_bot_64x8m81_0/nmos_5p04310589983270_64x8m81_0/D pmos_5p04310589983273_64x8m81_0/D
+ vdd xpredec0_bot_64x8m81_0/pmos_1p2$$47504428_64x8m81_0/pmos_5p04310589983267_64x8m81_0/D
+ xpredec0_bot_64x8m81_0/nmos_5p04310589983270_64x8m81_0/D xpredec0_bot_64x8m81_1/pmos_1p2$$47504428_64x8m81_0/pmos_5p04310589983267_64x8m81_0/D
+ A[0] vdd xpredec0_bot_64x8m81_1/nmos_5p04310589983270_64x8m81_0/D vss nmos_5p04310589983240_64x8m81_1/S
+ xpredec0_bot_64x8m81
Xxpredec0_bot_64x8m81_1 xpredec0_bot_64x8m81_0/pmos_1p2$$47504428_64x8m81_0/pmos_5p04310589983267_64x8m81_0/D
+ xpredec0_bot_64x8m81_0/nmos_5p04310589983270_64x8m81_0/D pmos_5p04310589983273_64x8m81_0/D
+ vdd xpredec0_bot_64x8m81_1/pmos_1p2$$47504428_64x8m81_0/pmos_5p04310589983267_64x8m81_0/D
+ xpredec0_bot_64x8m81_1/nmos_5p04310589983270_64x8m81_0/D xpredec0_bot_64x8m81_1/pmos_1p2$$47504428_64x8m81_0/pmos_5p04310589983267_64x8m81_0/D
+ A[1] vdd xpredec0_bot_64x8m81_1/nmos_5p04310589983270_64x8m81_0/D vss nmos_5p04310589983240_64x8m81_1/S
+ xpredec0_bot_64x8m81
Xpmos_5p04310589983273_64x8m81_0 vdd pmos_5p04310589983273_64x8m81_0/D nmos_5p04310589983240_64x8m81_1/S
+ vdd nmos_5p04310589983240_64x8m81_1/S pmos_5p04310589983273_64x8m81
Xnmos_5p04310589983240_64x8m81_0 nmos_5p04310589983240_64x8m81_1/S men vss vss nmos_5p04310589983240_64x8m81
Xnmos_5p04310589983240_64x8m81_1 vss clk nmos_5p04310589983240_64x8m81_1/S vss nmos_5p04310589983240_64x8m81
Xxpredec0_xa_64x8m81_0 xpredec0_xa_64x8m81_2/nmos_1p2$$47641644_64x8m81_0/nmos_5p04310589983261_64x8m81_0/S
+ xpredec0_bot_64x8m81_0/nmos_5p04310589983270_64x8m81_0/D xpredec0_bot_64x8m81_0/pmos_1p2$$47504428_64x8m81_0/pmos_5p04310589983267_64x8m81_0/D
+ vdd xpredec0_bot_64x8m81_1/pmos_1p2$$47504428_64x8m81_0/pmos_5p04310589983267_64x8m81_0/D
+ xpredec0_bot_64x8m81_1/pmos_1p2$$47504428_64x8m81_0/pmos_5p04310589983267_64x8m81_0/D
+ vss x[0] xpredec0_bot_64x8m81_0/pmos_1p2$$47504428_64x8m81_0/pmos_5p04310589983267_64x8m81_0/D
+ xpredec0_bot_64x8m81_1/nmos_5p04310589983270_64x8m81_0/D vdd vss vss vdd xpredec0_xa_64x8m81
Xxpredec0_xa_64x8m81_2 xpredec0_xa_64x8m81_2/nmos_1p2$$47641644_64x8m81_0/nmos_5p04310589983261_64x8m81_0/S
+ xpredec0_bot_64x8m81_0/nmos_5p04310589983270_64x8m81_0/D xpredec0_bot_64x8m81_0/nmos_5p04310589983270_64x8m81_0/D
+ vdd xpredec0_bot_64x8m81_1/pmos_1p2$$47504428_64x8m81_0/pmos_5p04310589983267_64x8m81_0/D
+ xpredec0_bot_64x8m81_1/pmos_1p2$$47504428_64x8m81_0/pmos_5p04310589983267_64x8m81_0/D
+ vss x[1] xpredec0_bot_64x8m81_0/pmos_1p2$$47504428_64x8m81_0/pmos_5p04310589983267_64x8m81_0/D
+ xpredec0_bot_64x8m81_1/nmos_5p04310589983270_64x8m81_0/D vdd vss vss vdd xpredec0_xa_64x8m81
Xxpredec0_xa_64x8m81_1 xpredec0_xa_64x8m81_3/nmos_1p2$$47641644_64x8m81_0/nmos_5p04310589983261_64x8m81_0/S
+ xpredec0_bot_64x8m81_0/nmos_5p04310589983270_64x8m81_0/D xpredec0_bot_64x8m81_0/pmos_1p2$$47504428_64x8m81_0/pmos_5p04310589983267_64x8m81_0/D
+ vdd xpredec0_bot_64x8m81_1/nmos_5p04310589983270_64x8m81_0/D xpredec0_bot_64x8m81_1/pmos_1p2$$47504428_64x8m81_0/pmos_5p04310589983267_64x8m81_0/D
+ vss x[2] xpredec0_bot_64x8m81_0/pmos_1p2$$47504428_64x8m81_0/pmos_5p04310589983267_64x8m81_0/D
+ xpredec0_bot_64x8m81_1/nmos_5p04310589983270_64x8m81_0/D vdd vss vss vdd xpredec0_xa_64x8m81
Xxpredec0_xa_64x8m81_3 xpredec0_xa_64x8m81_3/nmos_1p2$$47641644_64x8m81_0/nmos_5p04310589983261_64x8m81_0/S
+ xpredec0_bot_64x8m81_0/nmos_5p04310589983270_64x8m81_0/D xpredec0_bot_64x8m81_0/nmos_5p04310589983270_64x8m81_0/D
+ vdd xpredec0_bot_64x8m81_1/nmos_5p04310589983270_64x8m81_0/D xpredec0_bot_64x8m81_1/pmos_1p2$$47504428_64x8m81_0/pmos_5p04310589983267_64x8m81_0/D
+ vss x[3] xpredec0_bot_64x8m81_0/pmos_1p2$$47504428_64x8m81_0/pmos_5p04310589983267_64x8m81_0/D
+ xpredec0_bot_64x8m81_1/nmos_5p04310589983270_64x8m81_0/D vdd vss vss vdd xpredec0_xa_64x8m81
Xnmos_1p2$$46563372_64x8m81_0 pmos_5p04310589983273_64x8m81_0/D vss nmos_5p04310589983240_64x8m81_1/S
+ vss nmos_1p2$$46563372_64x8m81
X0 vdd men a_4894_9505# vdd pmos_3p3 w=1.705u l=0.6u
X1 a_4446_9505# men vdd vdd pmos_3p3 w=1.705u l=0.6u
X2 a_4894_9505# clk nmos_5p04310589983240_64x8m81_1/S vdd pmos_3p3 w=1.705u l=0.6u
X3 nmos_5p04310589983240_64x8m81_1/S clk a_4446_9505# vdd pmos_3p3 w=1.705u l=0.6u
.ends

.subckt prexdec_top_64x8m81 clk A[2] A[6] A[4] xb[3] xa[0] xc[0] xc[1] xc[2] xc[3]
+ xb[1] xb[2] xb[0] xa[1] xa[2] xa[3] xa[4] xa[5] xa[6] xa[7] A[0] A[3] A[5] A[1]
+ xpredec0_64x8m81_1/xpredec0_xa_64x8m81_2/nmos_1p2$$47641644_64x8m81_0/nmos_5p04310589983261_64x8m81_0/S
+ xpredec0_64x8m81_1/xpredec0_xa_64x8m81_3/nmos_1p2$$47641644_64x8m81_0/nmos_5p04310589983261_64x8m81_0/S
+ xpredec0_64x8m81_0/xpredec0_xa_64x8m81_2/nmos_1p2$$47641644_64x8m81_0/nmos_5p04310589983261_64x8m81_0/S
+ xpredec0_64x8m81_0/xpredec0_xa_64x8m81_3/nmos_1p2$$47641644_64x8m81_0/nmos_5p04310589983261_64x8m81_0/S
+ xpredec1_64x8m81_0/pmos_1p2$$47109164_64x8m81_0/pmos_5p04310589983266_64x8m81_0/w_n208_n120#
+ xpredec1_64x8m81_0/w_7178_9364# men xpredec1_64x8m81_0/vdd VSUBS
Xxpredec1_64x8m81_0 A[2] men xa[7] xa[6] xa[5] xa[4] xa[3] xa[2] xa[1] xa[0] A[1]
+ A[0] clk xpredec1_64x8m81_0/w_7178_9364# xpredec1_64x8m81_0/vdd xpredec1_64x8m81_0/pmos_1p2$$47109164_64x8m81_0/pmos_5p04310589983266_64x8m81_0/w_n208_n120#
+ VSUBS xpredec1_64x8m81
Xxpredec0_64x8m81_1 A[5] men xc[0] xc[1] xc[2] xc[3] A[6] clk xpredec0_64x8m81_1/xpredec0_xa_64x8m81_2/nmos_1p2$$47641644_64x8m81_0/nmos_5p04310589983261_64x8m81_0/S
+ xpredec0_64x8m81_1/xpredec0_xa_64x8m81_3/nmos_1p2$$47641644_64x8m81_0/nmos_5p04310589983261_64x8m81_0/S
+ VSUBS xpredec1_64x8m81_0/vdd xpredec0_64x8m81
Xxpredec0_64x8m81_0 A[3] men xb[0] xb[1] xb[2] xb[3] A[4] clk xpredec0_64x8m81_0/xpredec0_xa_64x8m81_2/nmos_1p2$$47641644_64x8m81_0/nmos_5p04310589983261_64x8m81_0/S
+ xpredec0_64x8m81_0/xpredec0_xa_64x8m81_3/nmos_1p2$$47641644_64x8m81_0/nmos_5p04310589983261_64x8m81_0/S
+ VSUBS xpredec1_64x8m81_0/vdd xpredec0_64x8m81
.ends

.subckt control_512x8_64x8m81 GWE GWEN VSS VDD RYS[7] RYS[6] RYS[5] RYS[4] RYS[3]
+ RYS[1] RYS[0] LYS[0] LYS[1] LYS[2] LYS[3] LYS[6] LYS[5] LYS[4] LYS[7] tblhl xb[3]
+ xb[2] xb[0] xa[7] xa[5] xa[4] xa[3] xa[2] A[0] xb[1] xc[3] xc[1] xc[2] xc[0] xa[0]
+ xa[1] A[9] A[7] CLK A[2] A[1] A[6] A[3] A[4] A[5] A[8] ypredec1_64x8m81_0/ly[2]
+ gen_512x8_64x8m81_0/tblhl IGWEN gen_512x8_64x8m81_0/wen_v2_64x8m81_0/nmos_5p0431058998329_64x8m81_4/D
+ CEN xa[6] RYS[2] ypredec1_64x8m81_0/ypredec1_bot_64x8m81_2/alatch_64x8m81_0/vdd
+ men prexdec_top_64x8m81_0/xpredec1_64x8m81_0/vdd VSUBS gen_512x8_64x8m81_0/VDD
Xgen_512x8_64x8m81_0 GWEN GWE gen_512x8_64x8m81_0/tblhl CEN CLK IGWEN gen_512x8_64x8m81_0/pmos_5p04310589983292_64x8m81_0/D
+ gen_512x8_64x8m81_0/wen_v2_64x8m81_0/nmos_5p0431058998329_64x8m81_4/D men VSUBS
+ gen_512x8_64x8m81_0/VDD gen_512x8_64x8m81
Xypredec1_64x8m81_0 ypredec1_64x8m81_0/ly[5] ypredec1_64x8m81_0/ly[4] ypredec1_64x8m81_0/ly[7]
+ ypredec1_64x8m81_0/ly[3] ypredec1_64x8m81_0/ly[2] ypredec1_64x8m81_0/ly[1] ypredec1_64x8m81_0/ly[0]
+ RYS[0] RYS[1] RYS[2] RYS[3] RYS[4] RYS[5] RYS[6] RYS[7] ypredec1_64x8m81_0/ly[6]
+ men A[0] A[1] A[2] CLK gen_512x8_64x8m81_0/VDD ypredec1_64x8m81_0/ypredec1_bot_64x8m81_2/alatch_64x8m81_0/vdd
+ VSUBS gen_512x8_64x8m81_0/VDD gen_512x8_64x8m81_0/VDD gen_512x8_64x8m81_0/VDD ypredec1_64x8m81
Xprexdec_top_64x8m81_0 CLK A[5] A[9] A[7] xb[3] xa[0] xc[0] xc[1] xc[2] xc[3] xb[1]
+ xb[2] xb[0] xa[1] xa[2] xa[3] xa[4] xa[5] xa[6] xa[7] A[3] A[6] A[8] A[4] VSUBS
+ VSUBS VSUBS VSUBS prexdec_top_64x8m81_0/xpredec1_64x8m81_0/vdd prexdec_top_64x8m81_0/xpredec1_64x8m81_0/vdd
+ men prexdec_top_64x8m81_0/xpredec1_64x8m81_0/vdd VSUBS prexdec_top_64x8m81
.ends

.subckt dcap_103_novia_64x8m81 w_n203_44# a_n67_185# a_73_103#
X0 a_n67_185# a_73_103# a_n67_185# w_n203_44# pmos_3p3 w=2.275u l=2.365u
.ends

.subckt pmos_5p04310589983218_64x8m81 w_n208_n120# D a_0_n44# a_896_n44# a_672_n44#
+ S a_448_n44# a_224_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X5 S a_1120_n44# D w_n208_n120# pmos_6p0 w=2.27u l=0.6u
.ends

.subckt pmos_1p2$$46549036_64x8m81 pmos_5p04310589983218_64x8m81_0/S a_193_n74# w_n286_n142#
+ a_1089_n74# a_865_n74# a_n31_n74# a_641_n74# pmos_5p04310589983218_64x8m81_0/D a_417_n74#
Xpmos_5p04310589983218_64x8m81_0 w_n286_n142# pmos_5p04310589983218_64x8m81_0/D a_n31_n74#
+ a_865_n74# a_641_n74# pmos_5p04310589983218_64x8m81_0/S a_417_n74# a_193_n74# a_1089_n74#
+ pmos_5p04310589983218_64x8m81
.ends

.subckt pmos_5p04310589983221_64x8m81 w_n208_n120# D a_0_n44# a_672_n44# S a_448_n44#
+ a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=0.91u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=0.91u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=0.91u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=0.91u l=0.6u
.ends

.subckt pmos_1p2$$46896172_64x8m81 pmos_5p04310589983221_64x8m81_0/S pmos_5p04310589983221_64x8m81_0/D
+ w_n286_n142# a_668_n74# a_n31_n74# a_193_n74# a_417_n74#
Xpmos_5p04310589983221_64x8m81_0 w_n286_n142# pmos_5p04310589983221_64x8m81_0/D a_n31_n74#
+ a_668_n74# pmos_5p04310589983221_64x8m81_0/S a_417_n74# a_193_n74# pmos_5p04310589983221_64x8m81
.ends

.subckt nmos_5p04310589983216_64x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# a_1568_n44# a_1344_n44# a_1120_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=3.41u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=3.41u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=3.41u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=3.41u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=3.41u l=0.6u
X5 S a_1120_n44# D VSUBS nmos_6p0 w=3.41u l=0.6u
X6 D a_1344_n44# S VSUBS nmos_6p0 w=3.41u l=0.6u
X7 S a_1568_n44# D VSUBS nmos_6p0 w=3.41u l=0.6u
.ends

.subckt nmos_1p2$$46552108_64x8m81 a_1089_n74# a_865_n74# a_641_n74# a_n31_n74# nmos_5p04310589983216_64x8m81_0/D
+ a_417_n74# a_193_n74# a_1537_n74# a_1313_n74# nmos_5p04310589983216_64x8m81_0/S
+ VSUBS
Xnmos_5p04310589983216_64x8m81_0 nmos_5p04310589983216_64x8m81_0/D a_n31_n74# a_865_n74#
+ a_641_n74# nmos_5p04310589983216_64x8m81_0/S a_417_n74# a_193_n74# a_1537_n74# a_1313_n74#
+ a_1089_n74# VSUBS nmos_5p04310589983216_64x8m81
.ends

.subckt nmos_5p04310589983217_64x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# a_1568_n44# a_1344_n44# a_1120_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.84u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2.84u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2.84u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=2.84u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=2.84u l=0.6u
X5 S a_1120_n44# D VSUBS nmos_6p0 w=2.84u l=0.6u
X6 D a_1344_n44# S VSUBS nmos_6p0 w=2.84u l=0.6u
X7 S a_1568_n44# D VSUBS nmos_6p0 w=2.84u l=0.6u
.ends

.subckt nmos_1p2$$46550060_64x8m81 a_1537_n74# a_1313_n74# nmos_5p04310589983217_64x8m81_0/D
+ a_193_n74# a_1089_n74# a_865_n74# a_n31_n74# a_641_n74# a_417_n74# VSUBS nmos_5p04310589983217_64x8m81_0/S
Xnmos_5p04310589983217_64x8m81_0 nmos_5p04310589983217_64x8m81_0/D a_n31_n74# a_865_n74#
+ a_641_n74# nmos_5p04310589983217_64x8m81_0/S a_417_n74# a_193_n74# a_1537_n74# a_1313_n74#
+ a_1089_n74# VSUBS nmos_5p04310589983217_64x8m81
.ends

.subckt pmos_1p2$$46897196_64x8m81 pmos_5p04310589983220_64x8m81_0/S pmos_5p04310589983220_64x8m81_0/D
+ a_193_n74# w_n286_n142# a_n31_n74#
Xpmos_5p04310589983220_64x8m81_0 w_n286_n142# pmos_5p04310589983220_64x8m81_0/D a_n31_n74#
+ pmos_5p04310589983220_64x8m81_0/S a_193_n74# pmos_5p04310589983220_64x8m81
.ends

.subckt pmos_5p04310589983219_64x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=0.91u l=0.6u
.ends

.subckt pmos_1p2$$46898220_64x8m81 pmos_5p04310589983219_64x8m81_0/S w_n286_n142#
+ a_n31_n74# pmos_5p04310589983219_64x8m81_0/D
Xpmos_5p04310589983219_64x8m81_0 w_n286_n142# pmos_5p04310589983219_64x8m81_0/D a_n31_n74#
+ pmos_5p04310589983219_64x8m81_0/S pmos_5p04310589983219_64x8m81
.ends

.subckt nmos_5p04310589983212_64x8m81 D a_0_n44# a_672_n44# S a_448_n44# a_224_n44#
+ VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
.ends

.subckt nmos_1p2$$45107244_64x8m81 a_193_n73# nmos_5p04310589983212_64x8m81_0/D a_n31_n73#
+ a_641_n73# a_417_n73# nmos_5p04310589983212_64x8m81_0/S VSUBS
Xnmos_5p04310589983212_64x8m81_0 nmos_5p04310589983212_64x8m81_0/D a_n31_n73# a_641_n73#
+ nmos_5p04310589983212_64x8m81_0/S a_417_n73# a_193_n73# VSUBS nmos_5p04310589983212_64x8m81
.ends

.subckt nmos_5p04310589983215_64x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=3.41u l=0.6u
.ends

.subckt nmos_1p2$$46553132_64x8m81 nmos_5p04310589983215_64x8m81_0/D a_n31_n74# nmos_5p04310589983215_64x8m81_0/S
+ VSUBS
Xnmos_5p04310589983215_64x8m81_0 nmos_5p04310589983215_64x8m81_0/D a_n31_n74# nmos_5p04310589983215_64x8m81_0/S
+ VSUBS nmos_5p04310589983215_64x8m81
.ends

.subckt pmos_5p04310589983213_64x8m81 w_n208_n120# D a_0_n44# S a_448_n44# a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
.ends

.subckt pmos_1p2$$46286892_64x8m81 a_193_n73# pmos_5p04310589983213_64x8m81_0/S a_n31_n73#
+ a_417_n73# w_n286_n142# pmos_5p04310589983213_64x8m81_0/D
Xpmos_5p04310589983213_64x8m81_0 w_n286_n142# pmos_5p04310589983213_64x8m81_0/D a_n31_n73#
+ pmos_5p04310589983213_64x8m81_0/S a_417_n73# a_193_n73# pmos_5p04310589983213_64x8m81
.ends

.subckt sa_64x8m81 wep se pcb qp d vss
Xpmos_1p2$$46549036_64x8m81_0 d pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S
+ d pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S
+ pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S qp qp qp pmos_1p2$$46549036_64x8m81
Xpmos_1p2$$46896172_64x8m81_0 pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S
+ d d pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S
+ pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S
+ pmos_1p2$$46896172_64x8m81
Xnmos_1p2$$46552108_64x8m81_0 pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S
+ pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S
+ pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S nmos_1p2$$46552108_64x8m81_0/nmos_5p04310589983216_64x8m81_0/D
+ pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S
+ pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S
+ pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S vss nmos_1p2$$46552108_64x8m81
Xnmos_1p2$$46550060_64x8m81_0 se se nmos_1p2$$46552108_64x8m81_0/nmos_5p04310589983216_64x8m81_0/D
+ se se se se se se vss vss nmos_1p2$$46550060_64x8m81
Xpmos_1p2$$46897196_64x8m81_0 d pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S
+ se d se pmos_1p2$$46897196_64x8m81
Xpmos_1p2$$46897196_64x8m81_1 d pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S
+ se d se pmos_1p2$$46897196_64x8m81
Xnmos_1p2$$46551084_64x8m81_0 vss pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S
+ qp vss nmos_1p2$$46551084_64x8m81
Xpmos_1p2$$46897196_64x8m81_2 d pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S
+ se d se pmos_1p2$$46897196_64x8m81
Xpmos_1p2$$46897196_64x8m81_3 d pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S
+ se d se pmos_1p2$$46897196_64x8m81
Xpmos_1p2$$46285868_64x8m81_0 pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S
+ d pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S pcb pmos_1p2$$46285868_64x8m81
Xpmos_1p2$$46898220_64x8m81_0 d d d pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S
+ pmos_1p2$$46898220_64x8m81
Xnmos_1p2$$45107244_64x8m81_0 qp vss pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S
+ qp qp qp vss nmos_1p2$$45107244_64x8m81
Xpmos_1p2$$46898220_64x8m81_1 pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S
+ d d d pmos_1p2$$46898220_64x8m81
Xnmos_1p2$$46553132_64x8m81_0 vss vss pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S
+ vss nmos_1p2$$46553132_64x8m81
Xnmos_1p2$$46553132_64x8m81_1 pmos_1p2$$46898220_64x8m81_1/pmos_5p04310589983219_64x8m81_0/S
+ vss vss vss nmos_1p2$$46553132_64x8m81
Xpmos_1p2$$46286892_64x8m81_0 pcb d pcb pcb d d pmos_1p2$$46286892_64x8m81
.ends

.subckt pmos_1p2$$202585132_64x8m81 w_n256_n141# pmos_5p04310589983214_64x8m81_0/S
+ pmos_5p04310589983214_64x8m81_0/D a_n31_n74#
Xpmos_5p04310589983214_64x8m81_0 w_n256_n141# pmos_5p04310589983214_64x8m81_0/D a_n31_n74#
+ pmos_5p04310589983214_64x8m81_0/S pmos_5p04310589983214_64x8m81
.ends

.subckt nmos_1p2$$202598444_64x8m81 nmos_5p0431058998325_64x8m81_0/D a_n31_n74# nmos_5p0431058998325_64x8m81_0/S
+ VSUBS
Xnmos_5p0431058998325_64x8m81_0 nmos_5p0431058998325_64x8m81_0/D a_n31_n74# nmos_5p0431058998325_64x8m81_0/S
+ VSUBS nmos_5p0431058998325_64x8m81
.ends

.subckt pmos_5p04310589983234_64x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=1.71u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.71u l=0.6u
.ends

.subckt nmos_1p2$$202594348_64x8m81 a_n31_n73# nmos_5p04310589983240_64x8m81_0/S nmos_5p04310589983240_64x8m81_0/D
+ VSUBS
Xnmos_5p04310589983240_64x8m81_0 nmos_5p04310589983240_64x8m81_0/D a_n31_n73# nmos_5p04310589983240_64x8m81_0/S
+ VSUBS nmos_5p04310589983240_64x8m81
.ends

.subckt pmos_1p2$$202584108_64x8m81 pmos_5p04310589983214_64x8m81_0/S a_n31_n74# w_n286_n141#
+ pmos_5p04310589983214_64x8m81_0/D
Xpmos_5p04310589983214_64x8m81_0 w_n286_n141# pmos_5p04310589983214_64x8m81_0/D a_n31_n74#
+ pmos_5p04310589983214_64x8m81_0/S pmos_5p04310589983214_64x8m81
.ends

.subckt pmos_5p04310589983242_64x8m81 w_n208_n120# D a_0_n44# S a_448_n44# a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=2u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=2u l=0.6u
.ends

.subckt pmos_1p2$$202583084_64x8m81 pmos_5p04310589983234_64x8m81_0/D a_193_n74# w_n286_n142#
+ a_n31_n74# pmos_5p04310589983234_64x8m81_0/S
Xpmos_5p04310589983234_64x8m81_0 w_n286_n142# pmos_5p04310589983234_64x8m81_0/D a_n31_n74#
+ pmos_5p04310589983234_64x8m81_0/S a_193_n74# pmos_5p04310589983234_64x8m81
.ends

.subckt nmos_5p04310589983243_64x8m81 D a_0_n44# S a_448_n44# a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=0.8u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=0.8u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=0.8u l=0.6u
.ends

.subckt wen_wm1_64x8m81 wep wen GWEN vss men vdd
Xnmos_1p2$$202596396_64x8m81_1 pmos_5p04310589983241_64x8m81_0/D vss nmos_1p2$$202595372_64x8m81_1/nmos_5p0431058998329_64x8m81_0/S
+ vss nmos_1p2$$202596396_64x8m81
Xnmos_5p0431058998329_64x8m81_3 nmos_5p0431058998329_64x8m81_3/D pmos_5p04310589983214_64x8m81_5/D
+ vss vss nmos_5p0431058998329_64x8m81
Xpmos_1p2$$202585132_64x8m81_0 vdd vdd nmos_1p2$$202596396_64x8m81_0/nmos_5p0431058998329_64x8m81_0/D
+ nmos_1p2$$202595372_64x8m81_1/nmos_5p0431058998329_64x8m81_0/S pmos_1p2$$202585132_64x8m81
Xpmos_1p2$$202586156_64x8m81_0 pmos_5p04310589983241_64x8m81_0/D vdd vdd nmos_1p2$$202595372_64x8m81_1/nmos_5p0431058998329_64x8m81_0/S
+ pmos_1p2$$202586156_64x8m81
Xnmos_1p2$$202598444_64x8m81_0 pmos_5p04310589983241_64x8m81_0/S pmos_5p04310589983214_64x8m81_5/D
+ nmos_5p0431058998329_64x8m81_1/D vss nmos_1p2$$202598444_64x8m81
Xpmos_5p04310589983234_64x8m81_0 vdd pmos_5p04310589983234_64x8m81_0/D nmos_5p0431058998325_64x8m81_0/S
+ vdd nmos_5p0431058998325_64x8m81_0/S pmos_5p04310589983234_64x8m81
Xnmos_5p04310589983239_64x8m81_0 men pmos_1p2$$202583084_64x8m81_0/pmos_5p04310589983234_64x8m81_0/D
+ nmos_5p0431058998325_64x8m81_0/S pmos_1p2$$202583084_64x8m81_0/pmos_5p04310589983234_64x8m81_0/D
+ vss nmos_5p04310589983239_64x8m81
Xpmos_5p04310589983220_64x8m81_0 vdd men nmos_1p2$$202596396_64x8m81_0/nmos_5p0431058998329_64x8m81_0/D
+ nmos_5p0431058998325_64x8m81_0/S nmos_1p2$$202596396_64x8m81_0/nmos_5p0431058998329_64x8m81_0/D
+ pmos_5p04310589983220_64x8m81
Xnmos_5p04310589983240_64x8m81_0 pmos_5p04310589983234_64x8m81_0/D nmos_5p0431058998325_64x8m81_0/S
+ vss vss nmos_5p04310589983240_64x8m81
Xpmos_1p2$$202587180_64x8m81_0 nmos_5p0431058998329_64x8m81_1/D vdd pmos_5p04310589983241_64x8m81_0/S
+ nmos_5p0431058998329_64x8m81_3/D pmos_1p2$$202587180_64x8m81
Xnmos_5p04310589983240_64x8m81_1 pmos_5p04310589983214_64x8m81_5/D men vss vss nmos_5p04310589983240_64x8m81
Xpmos_5p04310589983214_64x8m81_0 vdd pmos_5p04310589983214_64x8m81_2/S wen vdd pmos_5p04310589983214_64x8m81
Xnmos_5p04310589983240_64x8m81_2 vss vss pmos_5p04310589983214_64x8m81_5/D vss nmos_5p04310589983240_64x8m81
Xnmos_1p2$$202594348_64x8m81_0 nmos_1p2$$202596396_64x8m81_0/nmos_5p0431058998329_64x8m81_0/D
+ pmos_1p2$$202583084_64x8m81_0/pmos_5p04310589983234_64x8m81_0/D vss vss nmos_1p2$$202594348_64x8m81
Xpmos_5p04310589983214_64x8m81_1 vdd nmos_5p0431058998329_64x8m81_1/D nmos_5p0431058998329_64x8m81_2/D
+ vdd pmos_5p04310589983214_64x8m81
Xpmos_5p04310589983214_64x8m81_2 vdd nmos_5p0431058998329_64x8m81_2/D GWEN pmos_5p04310589983214_64x8m81_2/S
+ pmos_5p04310589983214_64x8m81
Xpmos_5p04310589983214_64x8m81_3 vdd pmos_5p04310589983214_64x8m81_5/S men vdd pmos_5p04310589983214_64x8m81
Xpmos_5p04310589983214_64x8m81_4 vdd nmos_5p0431058998329_64x8m81_3/D pmos_5p04310589983214_64x8m81_5/D
+ vdd pmos_5p04310589983214_64x8m81
Xpmos_5p04310589983214_64x8m81_5 vdd pmos_5p04310589983214_64x8m81_5/D vss pmos_5p04310589983214_64x8m81_5/S
+ pmos_5p04310589983214_64x8m81
Xpmos_1p2$$202584108_64x8m81_0 nmos_1p2$$202595372_64x8m81_1/nmos_5p0431058998329_64x8m81_0/S
+ pmos_5p04310589983241_64x8m81_0/S vdd vdd pmos_1p2$$202584108_64x8m81
Xpmos_5p04310589983242_64x8m81_0 vdd wep pmos_5p04310589983234_64x8m81_0/D vdd pmos_5p04310589983234_64x8m81_0/D
+ pmos_5p04310589983234_64x8m81_0/D pmos_5p04310589983242_64x8m81
Xpmos_1p2$$202583084_64x8m81_0 pmos_1p2$$202583084_64x8m81_0/pmos_5p04310589983234_64x8m81_0/D
+ nmos_1p2$$202596396_64x8m81_0/nmos_5p0431058998329_64x8m81_0/D vdd nmos_1p2$$202596396_64x8m81_0/nmos_5p0431058998329_64x8m81_0/D
+ vdd pmos_1p2$$202583084_64x8m81
Xnmos_5p04310589983243_64x8m81_0 wep pmos_5p04310589983234_64x8m81_0/D vss pmos_5p04310589983234_64x8m81_0/D
+ pmos_5p04310589983234_64x8m81_0/D vss nmos_5p04310589983243_64x8m81
Xnmos_5p0431058998325_64x8m81_0 vss nmos_1p2$$202596396_64x8m81_0/nmos_5p0431058998329_64x8m81_0/D
+ nmos_5p0431058998325_64x8m81_0/S vss nmos_5p0431058998325_64x8m81
Xnmos_5p0431058998329_64x8m81_0 vss GWEN nmos_5p0431058998329_64x8m81_2/D vss nmos_5p0431058998329_64x8m81
Xnmos_1p2$$202595372_64x8m81_0 pmos_5p04310589983241_64x8m81_0/S pmos_5p04310589983241_64x8m81_0/D
+ nmos_5p0431058998329_64x8m81_3/D vss nmos_1p2$$202595372_64x8m81
Xnmos_1p2$$202595372_64x8m81_1 nmos_1p2$$202595372_64x8m81_1/nmos_5p0431058998329_64x8m81_0/S
+ vss pmos_5p04310589983241_64x8m81_0/S vss nmos_1p2$$202595372_64x8m81
Xnmos_5p0431058998329_64x8m81_1 nmos_5p0431058998329_64x8m81_1/D nmos_5p0431058998329_64x8m81_2/D
+ vss vss nmos_5p0431058998329_64x8m81
Xpmos_5p04310589983241_64x8m81_0 vdd pmos_5p04310589983241_64x8m81_0/D pmos_5p04310589983214_64x8m81_5/D
+ pmos_5p04310589983241_64x8m81_0/S pmos_5p04310589983241_64x8m81
Xnmos_1p2$$202596396_64x8m81_0 vss nmos_1p2$$202596396_64x8m81_0/nmos_5p0431058998329_64x8m81_0/D
+ nmos_1p2$$202595372_64x8m81_1/nmos_5p0431058998329_64x8m81_0/S vss nmos_1p2$$202596396_64x8m81
Xnmos_5p0431058998329_64x8m81_2 nmos_5p0431058998329_64x8m81_2/D wen vss vss nmos_5p0431058998329_64x8m81
.ends

.subckt pmos_5p04310589983226_64x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=1.2u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.2u l=0.6u
.ends

.subckt nmos_5p04310589983232_64x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=1.44u l=0.6u
.ends

.subckt pmos_5p04310589983224_64x8m81 w_n208_n120# D a_0_n44# S a_448_n44# a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=4.54u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=4.54u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=4.54u l=0.6u
.ends

.subckt pmos_1p2$$46281772_64x8m81 a_n31_n73# pmos_5p04310589983224_64x8m81_0/S pmos_5p04310589983224_64x8m81_0/D
+ w_n286_n142# a_193_n73# a_417_n73#
Xpmos_5p04310589983224_64x8m81_0 w_n286_n142# pmos_5p04310589983224_64x8m81_0/D a_n31_n73#
+ pmos_5p04310589983224_64x8m81_0/S a_417_n73# a_193_n73# pmos_5p04310589983224_64x8m81
.ends

.subckt pmos_5p04310589983223_64x8m81 w_n208_n120# D a_0_n44# a_896_n44# a_672_n44#
+ S a_448_n44# a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
.ends

.subckt pmos_1p2$$46282796_64x8m81 pmos_5p04310589983223_64x8m81_0/S a_193_n74# a_865_n74#
+ a_n31_n74# a_641_n74# pmos_5p04310589983223_64x8m81_0/D a_417_n74# w_n286_n142#
Xpmos_5p04310589983223_64x8m81_0 w_n286_n142# pmos_5p04310589983223_64x8m81_0/D a_n31_n74#
+ a_865_n74# a_641_n74# pmos_5p04310589983223_64x8m81_0/S a_417_n74# a_193_n74# pmos_5p04310589983223_64x8m81
.ends

.subckt pmos_5p04310589983229_64x8m81 w_n208_n120# D a_2016_n44# a_0_n44# a_896_n44#
+ a_672_n44# S a_1792_n44# a_448_n44# a_224_n44# a_1568_n44# a_1344_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X5 S a_2016_n44# D w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X6 S a_1120_n44# D w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X7 D a_1344_n44# S w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X8 S a_1568_n44# D w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X9 D a_1792_n44# S w_n208_n120# pmos_6p0 w=2.72u l=0.6u
.ends

.subckt pmos_1p2$$45095980_64x8m81 a_193_n74# pmos_5p04310589983229_64x8m81_0/S a_1089_n74#
+ a_865_n74# a_n31_n74# a_641_n74# a_1985_n74# a_1761_n74# a_417_n74# w_n286_n142#
+ pmos_5p04310589983229_64x8m81_0/D a_1537_n74# a_1313_n74#
Xpmos_5p04310589983229_64x8m81_0 w_n286_n142# pmos_5p04310589983229_64x8m81_0/D a_1985_n74#
+ a_n31_n74# a_865_n74# a_641_n74# pmos_5p04310589983229_64x8m81_0/S a_1761_n74# a_417_n74#
+ a_193_n74# a_1537_n74# a_1313_n74# a_1089_n74# pmos_5p04310589983229_64x8m81
.ends

.subckt nmos_5p04310589983231_64x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=1.14u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=1.14u l=0.6u
.ends

.subckt pmos_5p04310589983222_64x8m81 w_n208_n120# D a_2016_n44# a_0_n44# a_896_n44#
+ a_672_n44# S a_1792_n44# a_448_n44# a_224_n44# a_1568_n44# a_1344_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X5 S a_2016_n44# D w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X6 S a_1120_n44# D w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X7 D a_1344_n44# S w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X8 S a_1568_n44# D w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X9 D a_1792_n44# S w_n208_n120# pmos_6p0 w=4.09u l=0.6u
.ends

.subckt pmos_1p2$$46283820_64x8m81 a_641_n74# a_1985_n74# a_1761_n74# a_417_n74# pmos_5p04310589983222_64x8m81_0/S
+ a_1537_n74# a_1313_n74# pmos_5p04310589983222_64x8m81_0/D w_n286_n142# a_193_n74#
+ a_1089_n74# a_865_n74# a_n31_n74#
Xpmos_5p04310589983222_64x8m81_0 w_n286_n142# pmos_5p04310589983222_64x8m81_0/D a_1985_n74#
+ a_n31_n74# a_865_n74# a_641_n74# pmos_5p04310589983222_64x8m81_0/S a_1761_n74# a_417_n74#
+ a_193_n74# a_1537_n74# a_1313_n74# a_1089_n74# pmos_5p04310589983222_64x8m81
.ends

.subckt pmos_1p2$$46284844_64x8m81 a_n31_n74# pmos_5p04310589983234_64x8m81_0/D w_n286_n142#
+ a_193_n74# pmos_5p04310589983234_64x8m81_0/S
Xpmos_5p04310589983234_64x8m81_0 w_n286_n142# pmos_5p04310589983234_64x8m81_0/D a_n31_n74#
+ pmos_5p04310589983234_64x8m81_0/S a_193_n74# pmos_5p04310589983234_64x8m81
.ends

.subckt nmos_5p04310589983228_64x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.61u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=2.61u l=0.6u
.ends

.subckt nmos_1p2$$45100076_64x8m81 nmos_5p04310589983228_64x8m81_0/D a_193_n74# nmos_5p04310589983228_64x8m81_0/S
+ a_n31_n74# VSUBS
Xnmos_5p04310589983228_64x8m81_0 nmos_5p04310589983228_64x8m81_0/D a_n31_n74# nmos_5p04310589983228_64x8m81_0/S
+ a_193_n74# VSUBS nmos_5p04310589983228_64x8m81
.ends

.subckt pmos_5p04310589983233_64x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.2u l=0.6u
.ends

.subckt nmos_5p04310589983238_64x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=0.6u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=0.6u l=0.6u
.ends

.subckt nmos_5p04310589983235_64x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=1.14u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=1.14u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=1.14u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=1.14u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=1.14u l=0.6u
.ends

.subckt nmos_1p2$$45101100_64x8m81 a_193_n74# nmos_5p04310589983235_64x8m81_0/S a_865_n74#
+ a_n31_n74# a_641_n74# a_417_n74# nmos_5p04310589983235_64x8m81_0/D VSUBS
Xnmos_5p04310589983235_64x8m81_0 nmos_5p04310589983235_64x8m81_0/D a_n31_n74# a_865_n74#
+ a_641_n74# nmos_5p04310589983235_64x8m81_0/S a_417_n74# a_193_n74# VSUBS nmos_5p04310589983235_64x8m81
.ends

.subckt nmos_5p04310589983237_64x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=0.6u l=0.6u
.ends

.subckt nmos_5p04310589983225_64x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# a_1344_n44# a_1120_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X5 S a_1120_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X6 D a_1344_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
.ends

.subckt nmos_1p2$$45102124_64x8m81 a_1313_n74# nmos_5p04310589983225_64x8m81_0/D a_193_n74#
+ a_1089_n74# nmos_5p04310589983225_64x8m81_0/S a_865_n74# a_n31_n74# a_641_n74# a_417_n74#
+ VSUBS
Xnmos_5p04310589983225_64x8m81_0 nmos_5p04310589983225_64x8m81_0/D a_n31_n74# a_865_n74#
+ a_641_n74# nmos_5p04310589983225_64x8m81_0/S a_417_n74# a_193_n74# a_1313_n74# a_1089_n74#
+ VSUBS nmos_5p04310589983225_64x8m81
.ends

.subckt pmos_5p04310589983230_64x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=3.41u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=3.41u l=0.6u
.ends

.subckt pmos_1p2$$46287916_64x8m81 pmos_5p04310589983230_64x8m81_0/D a_193_n74# w_n286_n142#
+ a_n31_n74# pmos_5p04310589983230_64x8m81_0/S
Xpmos_5p04310589983230_64x8m81_0 w_n286_n142# pmos_5p04310589983230_64x8m81_0/D a_n31_n74#
+ pmos_5p04310589983230_64x8m81_0/S a_193_n74# pmos_5p04310589983230_64x8m81
.ends

.subckt nmos_5p04310589983236_64x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# a_1120_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.86u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2.86u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2.86u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=2.86u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=2.86u l=0.6u
X5 S a_1120_n44# D VSUBS nmos_6p0 w=2.86u l=0.6u
.ends

.subckt nmos_1p2$$45103148_64x8m81 a_865_n73# a_193_n74# nmos_5p04310589983236_64x8m81_0/S
+ a_1089_n74# a_n31_n74# a_641_n74# a_417_n74# nmos_5p04310589983236_64x8m81_0/D VSUBS
Xnmos_5p04310589983236_64x8m81_0 nmos_5p04310589983236_64x8m81_0/D a_n31_n74# a_865_n73#
+ a_641_n74# nmos_5p04310589983236_64x8m81_0/S a_417_n74# a_193_n74# a_1089_n74# VSUBS
+ nmos_5p04310589983236_64x8m81
.ends

.subckt nmos_5p04310589983227_64x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
.ends

.subckt sacntl_2_64x8m81 pcb se men pmos_1p2$$46282796_64x8m81_0/pmos_5p04310589983223_64x8m81_0/D
+ a_4718_983# nmos_5p04310589983238_64x8m81_1/D pmos_5p04310589983226_64x8m81_2/S
+ pmos_5p04310589983226_64x8m81_1/S a_4560_1922# a_2796_670# vdd vss
Xpmos_5p04310589983226_64x8m81_2 vdd vdd pmos_5p04310589983226_64x8m81_1/S pmos_5p04310589983226_64x8m81_2/S
+ pmos_5p04310589983226_64x8m81_2/S pmos_5p04310589983226_64x8m81
Xnmos_5p04310589983232_64x8m81_0 nmos_5p04310589983232_64x8m81_0/D pmos_5p04310589983226_64x8m81_1/S
+ vss vss nmos_5p04310589983232_64x8m81
Xpmos_1p2$$46281772_64x8m81_0 pmos_1p2$$46281772_64x8m81_1/pmos_5p04310589983224_64x8m81_0/S
+ pmos_1p2$$46281772_64x8m81_0/pmos_5p04310589983224_64x8m81_0/S vdd vdd pmos_1p2$$46281772_64x8m81_1/pmos_5p04310589983224_64x8m81_0/S
+ pmos_1p2$$46281772_64x8m81_1/pmos_5p04310589983224_64x8m81_0/S pmos_1p2$$46281772_64x8m81
Xpmos_1p2$$46281772_64x8m81_1 pmos_1p2$$46282796_64x8m81_0/pmos_5p04310589983223_64x8m81_0/D
+ pmos_1p2$$46281772_64x8m81_1/pmos_5p04310589983224_64x8m81_0/S vdd vdd nmos_5p04310589983232_64x8m81_0/D
+ nmos_5p04310589983227_64x8m81_1/S pmos_1p2$$46281772_64x8m81
Xpmos_1p2$$46282796_64x8m81_0 vdd men men men men pmos_1p2$$46282796_64x8m81_0/pmos_5p04310589983223_64x8m81_0/D
+ men vdd pmos_1p2$$46282796_64x8m81
Xnmos_5p04310589983212_64x8m81_0 se nmos_5p04310589983227_64x8m81_1/S nmos_5p04310589983227_64x8m81_1/S
+ vss nmos_5p04310589983227_64x8m81_1/S nmos_5p04310589983227_64x8m81_1/S vss nmos_5p04310589983212_64x8m81
Xpmos_1p2$$45095980_64x8m81_0 nmos_5p04310589983227_64x8m81_1/S vdd nmos_5p04310589983227_64x8m81_1/S
+ nmos_5p04310589983227_64x8m81_1/S nmos_5p04310589983227_64x8m81_1/S nmos_5p04310589983227_64x8m81_1/S
+ nmos_5p04310589983227_64x8m81_1/S nmos_5p04310589983227_64x8m81_1/S nmos_5p04310589983227_64x8m81_1/S
+ vdd se nmos_5p04310589983227_64x8m81_1/S nmos_5p04310589983227_64x8m81_1/S pmos_1p2$$45095980_64x8m81
Xnmos_5p04310589983231_64x8m81_0 nmos_5p04310589983231_64x8m81_0/D nmos_5p04310589983232_64x8m81_0/D
+ vss nmos_5p04310589983232_64x8m81_0/D vss nmos_5p04310589983231_64x8m81
Xpmos_1p2$$46283820_64x8m81_0 pmos_1p2$$46281772_64x8m81_0/pmos_5p04310589983224_64x8m81_0/S
+ pmos_1p2$$46281772_64x8m81_0/pmos_5p04310589983224_64x8m81_0/S pmos_1p2$$46281772_64x8m81_0/pmos_5p04310589983224_64x8m81_0/S
+ pmos_1p2$$46281772_64x8m81_0/pmos_5p04310589983224_64x8m81_0/S vdd pmos_1p2$$46281772_64x8m81_0/pmos_5p04310589983224_64x8m81_0/S
+ pmos_1p2$$46281772_64x8m81_0/pmos_5p04310589983224_64x8m81_0/S pcb vdd pmos_1p2$$46281772_64x8m81_0/pmos_5p04310589983224_64x8m81_0/S
+ pmos_1p2$$46281772_64x8m81_0/pmos_5p04310589983224_64x8m81_0/S pmos_1p2$$46281772_64x8m81_0/pmos_5p04310589983224_64x8m81_0/S
+ pmos_1p2$$46281772_64x8m81_0/pmos_5p04310589983224_64x8m81_0/S pmos_1p2$$46283820_64x8m81
Xpmos_1p2$$46284844_64x8m81_0 pmos_5p04310589983226_64x8m81_1/S nmos_5p04310589983232_64x8m81_0/D
+ vdd pmos_5p04310589983226_64x8m81_1/S vdd pmos_1p2$$46284844_64x8m81
Xnmos_1p2$$45100076_64x8m81_0 pmos_1p2$$46281772_64x8m81_0/pmos_5p04310589983224_64x8m81_0/S
+ pmos_1p2$$46281772_64x8m81_1/pmos_5p04310589983224_64x8m81_0/S vss pmos_1p2$$46281772_64x8m81_1/pmos_5p04310589983224_64x8m81_0/S
+ vss nmos_1p2$$45100076_64x8m81
Xpmos_1p2$$46285868_64x8m81_0 nmos_5p04310589983227_64x8m81_1/S vdd vdd pmos_1p2$$46282796_64x8m81_0/pmos_5p04310589983223_64x8m81_0/D
+ pmos_1p2$$46285868_64x8m81
Xpmos_5p04310589983233_64x8m81_0 vdd vdd pmos_5p04310589983226_64x8m81_0/S pmos_5p04310589983233_64x8m81_0/S
+ pmos_5p04310589983233_64x8m81
Xnmos_5p04310589983238_64x8m81_0 vss a_2796_670# pmos_5p04310589983226_64x8m81_0/S
+ pmos_5p04310589983226_64x8m81_0/S vss nmos_5p04310589983238_64x8m81
Xnmos_5p04310589983238_64x8m81_1 nmos_5p04310589983238_64x8m81_1/D pmos_1p2$$46282796_64x8m81_0/pmos_5p04310589983223_64x8m81_0/D
+ pmos_5p04310589983226_64x8m81_1/S vss vss nmos_5p04310589983238_64x8m81
Xnmos_5p04310589983238_64x8m81_2 vss pmos_5p04310589983226_64x8m81_1/S pmos_5p04310589983226_64x8m81_2/S
+ pmos_5p04310589983226_64x8m81_2/S vss nmos_5p04310589983238_64x8m81
Xnmos_1p2$$45101100_64x8m81_0 men vss men men men men pmos_1p2$$46282796_64x8m81_0/pmos_5p04310589983223_64x8m81_0/D
+ vss nmos_1p2$$45101100_64x8m81
Xnmos_5p04310589983237_64x8m81_0 vss pmos_5p04310589983226_64x8m81_0/S pmos_5p04310589983233_64x8m81_0/S
+ vss nmos_5p04310589983237_64x8m81
Xnmos_1p2$$45102124_64x8m81_0 pmos_1p2$$46281772_64x8m81_0/pmos_5p04310589983224_64x8m81_0/S
+ pcb pmos_1p2$$46281772_64x8m81_0/pmos_5p04310589983224_64x8m81_0/S pmos_1p2$$46281772_64x8m81_0/pmos_5p04310589983224_64x8m81_0/S
+ vss pmos_1p2$$46281772_64x8m81_0/pmos_5p04310589983224_64x8m81_0/S pmos_1p2$$46281772_64x8m81_0/pmos_5p04310589983224_64x8m81_0/S
+ pmos_1p2$$46281772_64x8m81_0/pmos_5p04310589983224_64x8m81_0/S pmos_1p2$$46281772_64x8m81_0/pmos_5p04310589983224_64x8m81_0/S
+ vss nmos_1p2$$45102124_64x8m81
Xpmos_1p2$$46287916_64x8m81_0 nmos_5p04310589983231_64x8m81_0/D nmos_5p04310589983232_64x8m81_0/D
+ vdd nmos_5p04310589983232_64x8m81_0/D vdd pmos_1p2$$46287916_64x8m81
Xnmos_1p2$$45103148_64x8m81_0 nmos_5p04310589983232_64x8m81_0/D nmos_5p04310589983232_64x8m81_0/D
+ vss pmos_1p2$$46282796_64x8m81_0/pmos_5p04310589983223_64x8m81_0/D pmos_1p2$$46282796_64x8m81_0/pmos_5p04310589983223_64x8m81_0/D
+ nmos_5p04310589983227_64x8m81_1/S nmos_5p04310589983227_64x8m81_1/S pmos_1p2$$46281772_64x8m81_1/pmos_5p04310589983224_64x8m81_0/S
+ vss nmos_1p2$$45103148_64x8m81
Xpmos_5p04310589983226_64x8m81_0 vdd vdd a_2796_670# pmos_5p04310589983226_64x8m81_0/S
+ pmos_5p04310589983226_64x8m81_0/S pmos_5p04310589983226_64x8m81
Xnmos_5p04310589983227_64x8m81_0 nmos_5p04310589983227_64x8m81_1/D nmos_5p04310589983231_64x8m81_0/D
+ nmos_5p04310589983231_64x8m81_0/D nmos_5p04310589983231_64x8m81_0/D vss nmos_5p04310589983231_64x8m81_0/D
+ nmos_5p04310589983231_64x8m81_0/D vss nmos_5p04310589983227_64x8m81
Xpmos_1p2$$46286892_64x8m81_0 nmos_5p04310589983231_64x8m81_0/D vdd nmos_5p04310589983231_64x8m81_0/D
+ nmos_5p04310589983231_64x8m81_0/D vdd nmos_5p04310589983227_64x8m81_1/S pmos_1p2$$46286892_64x8m81
Xpmos_5p04310589983226_64x8m81_1 vdd vdd pmos_1p2$$46282796_64x8m81_0/pmos_5p04310589983223_64x8m81_0/D
+ pmos_5p04310589983226_64x8m81_1/S vss pmos_5p04310589983226_64x8m81
Xnmos_5p04310589983227_64x8m81_1 nmos_5p04310589983227_64x8m81_1/D pmos_1p2$$46282796_64x8m81_0/pmos_5p04310589983223_64x8m81_0/D
+ pmos_1p2$$46282796_64x8m81_0/pmos_5p04310589983223_64x8m81_0/D pmos_1p2$$46282796_64x8m81_0/pmos_5p04310589983223_64x8m81_0/D
+ nmos_5p04310589983227_64x8m81_1/S pmos_1p2$$46282796_64x8m81_0/pmos_5p04310589983223_64x8m81_0/D
+ pmos_1p2$$46282796_64x8m81_0/pmos_5p04310589983223_64x8m81_0/D vss nmos_5p04310589983227_64x8m81
.ends

.subckt nmos_5p04310589983245_64x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# a_1120_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.12u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2.12u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2.12u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=2.12u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=2.12u l=0.6u
X5 S a_1120_n44# D VSUBS nmos_6p0 w=2.12u l=0.6u
.ends

.subckt pmos_5p04310589983248_64x8m81 w_n208_n120# D a_0_n44# a_896_n44# a_672_n44#
+ S a_448_n44# a_224_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=3.78u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=3.78u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=3.78u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=3.78u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=3.78u l=0.6u
X5 S a_1120_n44# D w_n208_n120# pmos_6p0 w=3.78u l=0.6u
.ends

.subckt nmos_5p04310589983249_64x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=2.2u l=0.6u
.ends

.subckt pmos_1p2$$171625516_64x8m81 pmos_5p0431058998323_64x8m81_0/D a_193_n74# w_n286_n142#
+ pmos_5p0431058998323_64x8m81_0/w_n208_n120# pmos_5p0431058998323_64x8m81_0/S a_n31_n74#
Xpmos_5p0431058998323_64x8m81_0 pmos_5p0431058998323_64x8m81_0/w_n208_n120# pmos_5p0431058998323_64x8m81_0/D
+ a_n31_n74# pmos_5p0431058998323_64x8m81_0/S a_193_n74# pmos_5p0431058998323_64x8m81
.ends

.subckt nmos_5p04310589983250_64x8m81 D a_0_n44# S a_448_n44# a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
.ends

.subckt nmos_5p04310589983244_64x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.84u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=2.84u l=0.6u
.ends

.subckt pmos_5p04310589983247_64x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=4.5u l=0.6u
.ends

.subckt pmos_5p04310589983246_64x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=4u l=0.6u
.ends

.subckt nmos_5p04310589983252_64x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=1.6u l=0.6u
.ends

.subckt outbuf_oe_64x8m81 se q GWE qp qn a_4913_n316# vdd vss
Xnmos_5p04310589983245_64x8m81_0 vss pmos_5p04310589983251_64x8m81_0/D pmos_5p04310589983251_64x8m81_0/D
+ pmos_5p04310589983251_64x8m81_0/D q pmos_5p04310589983251_64x8m81_0/D pmos_5p04310589983251_64x8m81_0/D
+ pmos_5p04310589983251_64x8m81_0/D vss nmos_5p04310589983245_64x8m81
Xpmos_5p04310589983248_64x8m81_0 vdd vdd pmos_5p04310589983251_64x8m81_0/D pmos_5p04310589983251_64x8m81_0/D
+ pmos_5p04310589983251_64x8m81_0/D q pmos_5p04310589983251_64x8m81_0/D pmos_5p04310589983251_64x8m81_0/D
+ pmos_5p04310589983251_64x8m81_0/D pmos_5p04310589983248_64x8m81
Xnmos_5p04310589983249_64x8m81_0 vss pmos_5p04310589983246_64x8m81_0/S pmos_5p04310589983247_64x8m81_0/S
+ vss nmos_5p04310589983249_64x8m81
Xpmos_1p2$$171625516_64x8m81_0 nmos_5p0431058998329_64x8m81_1/S pmos_5p04310589983233_64x8m81_0/D
+ vdd vdd vdd pmos_5p04310589983233_64x8m81_0/D pmos_1p2$$171625516_64x8m81
Xnmos_5p04310589983250_64x8m81_0 nmos_5p0431058998329_64x8m81_1/S nmos_5p0431058998329_64x8m81_0/D
+ pmos_5p04310589983251_64x8m81_0/D nmos_5p0431058998329_64x8m81_0/D nmos_5p0431058998329_64x8m81_0/D
+ vss nmos_5p04310589983250_64x8m81
Xnmos_5p04310589983244_64x8m81_0 vss pmos_5p04310589983246_64x8m81_0/S nmos_5p04310589983244_64x8m81_1/S
+ pmos_5p04310589983246_64x8m81_0/S vss nmos_5p04310589983244_64x8m81
Xpmos_5p04310589983247_64x8m81_0 vdd vdd pmos_5p04310589983246_64x8m81_0/S pmos_5p04310589983247_64x8m81_0/S
+ pmos_5p04310589983247_64x8m81
Xpmos_5p04310589983214_64x8m81_0 vdd nmos_5p0431058998329_64x8m81_0/D se vdd pmos_5p04310589983214_64x8m81
Xnmos_5p04310589983244_64x8m81_1 pmos_5p04310589983251_64x8m81_0/D qn nmos_5p04310589983244_64x8m81_1/S
+ qn vss nmos_5p04310589983244_64x8m81
Xpmos_5p04310589983233_64x8m81_0 vdd pmos_5p04310589983233_64x8m81_0/D pmos_5p04310589983251_64x8m81_0/D
+ vdd pmos_5p04310589983233_64x8m81
Xpmos_5p04310589983213_64x8m81_0 vdd nmos_5p0431058998329_64x8m81_1/S se pmos_5p04310589983251_64x8m81_0/D
+ se se pmos_5p04310589983213_64x8m81
Xpmos_5p04310589983246_64x8m81_0 vdd vdd GWE pmos_5p04310589983246_64x8m81_0/S pmos_5p04310589983246_64x8m81
Xnmos_5p04310589983237_64x8m81_0 pmos_5p04310589983233_64x8m81_0/D pmos_5p04310589983251_64x8m81_0/D
+ vss vss nmos_5p04310589983237_64x8m81
Xpmos_5p04310589983251_64x8m81_0 vdd pmos_5p04310589983251_64x8m81_0/D qp pmos_5p04310589983251_64x8m81_1/S
+ qp pmos_5p04310589983251_64x8m81
Xpmos_5p04310589983251_64x8m81_1 vdd vdd pmos_5p04310589983247_64x8m81_0/S pmos_5p04310589983251_64x8m81_1/S
+ pmos_5p04310589983247_64x8m81_0/S pmos_5p04310589983251_64x8m81
Xnmos_5p04310589983252_64x8m81_0 vss GWE pmos_5p04310589983246_64x8m81_0/S vss nmos_5p04310589983252_64x8m81
Xnmos_5p0431058998329_64x8m81_0 nmos_5p0431058998329_64x8m81_0/D se vss vss nmos_5p0431058998329_64x8m81
Xnmos_5p0431058998329_64x8m81_1 vss pmos_5p04310589983233_64x8m81_0/D nmos_5p0431058998329_64x8m81_1/S
+ vss nmos_5p0431058998329_64x8m81
.ends

.subckt pmos_5p0431058998321_64x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=6.81u l=0.6u
.ends

.subckt pmos_1p2$$46889004_64x8m81 pmos_5p0431058998321_64x8m81_0/D w_n286_n142# pmos_5p0431058998321_64x8m81_0/S
+ a_n31_n74#
Xpmos_5p0431058998321_64x8m81_0 w_n286_n142# pmos_5p0431058998321_64x8m81_0/D a_n31_n74#
+ pmos_5p0431058998321_64x8m81_0/S pmos_5p0431058998321_64x8m81
.ends

.subckt pmos_5p04310589983210_64x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=11.34u l=0.6u
.ends

.subckt nmos_5p04310589983211_64x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=0.96u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=0.96u l=0.6u
.ends

.subckt pmos_5p0431058998327_64x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=0.96u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=0.96u l=0.6u
.ends

.subckt pmos_1p2$$46885932_64x8m81 a_193_n73# pmos_5p0431058998327_64x8m81_0/D a_n31_n74#
+ w_n286_n141# pmos_5p0431058998327_64x8m81_0/S
Xpmos_5p0431058998327_64x8m81_0 w_n286_n141# pmos_5p0431058998327_64x8m81_0/D a_n31_n74#
+ pmos_5p0431058998327_64x8m81_0/S a_193_n73# pmos_5p0431058998327_64x8m81
.ends

.subckt nmos_5p0431058998328_64x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=13.61u l=0.6u
.ends

.subckt nmos_1p2$$46884908_64x8m81 nmos_5p0431058998328_64x8m81_0/D a_n31_n74# VSUBS
+ nmos_5p0431058998328_64x8m81_0/S
Xnmos_5p0431058998328_64x8m81_0 nmos_5p0431058998328_64x8m81_0/D a_n31_n74# nmos_5p0431058998328_64x8m81_0/S
+ VSUBS nmos_5p0431058998328_64x8m81
.ends

.subckt nmos_5p0431058998326_64x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=11.34u l=0.6u
.ends

.subckt nmos_1p2$$46883884_64x8m81 nmos_5p0431058998326_64x8m81_0/D a_n31_n73# nmos_5p0431058998326_64x8m81_0/S
+ VSUBS
Xnmos_5p0431058998326_64x8m81_0 nmos_5p0431058998326_64x8m81_0/D a_n31_n73# nmos_5p0431058998326_64x8m81_0/S
+ VSUBS nmos_5p0431058998326_64x8m81
.ends

.subckt din_64x8m81 datain wep men d db pmos_5p0431058998321_64x8m81_0/D m1_164_8068#
+ vdd vss
Xnmos_1p2$$46563372_64x8m81_1 vss pmos_1p2$$46273580_64x8m81_0/pmos_5p0431058998323_64x8m81_0/D
+ men vss nmos_1p2$$46563372_64x8m81
Xpmos_1p2$$46887980_64x8m81_0 pmos_1p2$$46889004_64x8m81_0/pmos_5p0431058998321_64x8m81_0/D
+ vdd vdd pmos_5p0431058998321_64x8m81_0/S pmos_1p2$$46887980_64x8m81
Xpmos_5p0431058998321_64x8m81_0 vdd pmos_5p0431058998321_64x8m81_0/D nmos_5p04310589983211_64x8m81_1/D
+ pmos_5p0431058998321_64x8m81_0/S pmos_5p0431058998321_64x8m81
Xpmos_1p2$$46273580_64x8m81_0 pmos_1p2$$46273580_64x8m81_0/pmos_5p0431058998323_64x8m81_0/D
+ men vdd vdd men pmos_1p2$$46273580_64x8m81
Xpmos_1p2$$46273580_64x8m81_1 pmos_5p0431058998327_64x8m81_0/S pmos_5p0431058998321_64x8m81_0/S
+ vdd vdd pmos_5p0431058998321_64x8m81_0/S pmos_1p2$$46273580_64x8m81
Xpmos_1p2$$46889004_64x8m81_0 pmos_1p2$$46889004_64x8m81_0/pmos_5p0431058998321_64x8m81_0/D
+ vdd d a_500_6666# pmos_1p2$$46889004_64x8m81
Xpmos_5p04310589983210_64x8m81_0 vdd vdd pmos_1p2$$46889004_64x8m81_0/pmos_5p0431058998321_64x8m81_0/D
+ pmos_5p04310589983210_64x8m81_0/S pmos_5p04310589983210_64x8m81
Xnmos_5p04310589983211_64x8m81_0 vss datain pmos_5p0431058998327_64x8m81_0/S pmos_5p0431058998327_64x8m81_0/S
+ vss nmos_5p04310589983211_64x8m81
Xpmos_1p2$$46889004_64x8m81_1 pmos_5p04310589983210_64x8m81_0/S vdd db a_500_6666#
+ pmos_1p2$$46889004_64x8m81
Xnmos_5p04310589983211_64x8m81_1 nmos_5p04310589983211_64x8m81_1/D pmos_1p2$$46273580_64x8m81_0/pmos_5p0431058998323_64x8m81_0/D
+ pmos_5p0431058998327_64x8m81_0/S men vss nmos_5p04310589983211_64x8m81
Xpmos_1p2$$46885932_64x8m81_0 pmos_1p2$$46273580_64x8m81_0/pmos_5p0431058998323_64x8m81_0/D
+ nmos_5p04310589983211_64x8m81_1/D men vdd pmos_5p0431058998327_64x8m81_0/S pmos_1p2$$46885932_64x8m81
Xnmos_1p2$$46884908_64x8m81_0 pmos_1p2$$46889004_64x8m81_0/pmos_5p0431058998321_64x8m81_0/D
+ pmos_5p0431058998321_64x8m81_0/S vss vss nmos_1p2$$46884908_64x8m81
Xnmos_1p2$$46883884_64x8m81_0 pmos_5p04310589983210_64x8m81_0/S wep db vss nmos_1p2$$46883884_64x8m81
Xnmos_1p2$$46883884_64x8m81_1 vss pmos_1p2$$46889004_64x8m81_0/pmos_5p0431058998321_64x8m81_0/D
+ pmos_5p04310589983210_64x8m81_0/S vss nmos_1p2$$46883884_64x8m81
Xnmos_1p2$$46883884_64x8m81_2 pmos_1p2$$46889004_64x8m81_0/pmos_5p0431058998321_64x8m81_0/D
+ wep d vss nmos_1p2$$46883884_64x8m81
Xpmos_5p0431058998327_64x8m81_0 vdd vdd datain pmos_5p0431058998327_64x8m81_0/S pmos_5p0431058998327_64x8m81_0/S
+ pmos_5p0431058998327_64x8m81
Xnmos_5p0431058998325_64x8m81_0 vss nmos_5p04310589983211_64x8m81_1/D pmos_5p0431058998321_64x8m81_0/S
+ vss nmos_5p0431058998325_64x8m81
Xnmos_1p2$$46563372_64x8m81_0 vss pmos_5p0431058998327_64x8m81_0/S pmos_5p0431058998321_64x8m81_0/S
+ vss nmos_1p2$$46563372_64x8m81
X0 vdd wep a_500_6666# vdd pmos_3p3 w=1.485u l=0.6u
X1 a_500_6666# wep vss vss nmos_3p3 w=1.14u l=0.6u
X2 a_500_6666# wep vdd vdd pmos_3p3 w=1.485u l=0.6u
.ends

.subckt nmos_5p0431058998320_64x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=6.81u l=0.6u
.ends

.subckt nmos_1p2$$47119404_64x8m81 nmos_5p0431058998320_64x8m81_0/D nmos_5p0431058998320_64x8m81_0/S
+ a_n31_n74# VSUBS
Xnmos_5p0431058998320_64x8m81_0 nmos_5p0431058998320_64x8m81_0/D a_n31_n74# nmos_5p0431058998320_64x8m81_0/S
+ VSUBS nmos_5p0431058998320_64x8m81
.ends

.subckt nmos_5p0431058998322_64x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=0.57u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=0.57u l=0.6u
.ends

.subckt ypass_gate_a_64x8m81 d pcb vss b bb db ypass a_222_11191# a_n4_11191# m3_n1_4331#
+ a_447_11191# a_n80_n10# a_222_10416# m3_n1_1708# a_n4_10416# m3_n1_1160# m3_n1_2030#
+ vdd pmos_5p0431058998321_64x8m81_1/D m3_n1_3366# a_447_10416# m3_n1_2352# m3_n1_3688#
+ m3_n1_4009# m3_n1_2674#
Xpmos_5p0431058998321_64x8m81_0 vdd b pcb bb pmos_5p0431058998321_64x8m81
Xpmos_5p0431058998321_64x8m81_1 vdd pmos_5p0431058998321_64x8m81_1/D nmos_5p0431058998322_64x8m81_0/D
+ bb pmos_5p0431058998321_64x8m81
Xnmos_1p2$$47119404_64x8m81_0 d b ypass vss nmos_1p2$$47119404_64x8m81
Xnmos_1p2$$47119404_64x8m81_1 pmos_5p0431058998321_64x8m81_1/D bb ypass vss nmos_1p2$$47119404_64x8m81
Xpmos_1p2$$46889004_64x8m81_0 d vdd b nmos_5p0431058998322_64x8m81_0/D pmos_1p2$$46889004_64x8m81
Xnmos_5p0431058998322_64x8m81_0 nmos_5p0431058998322_64x8m81_0/D ypass vss ypass vss
+ nmos_5p0431058998322_64x8m81
X0 nmos_5p0431058998322_64x8m81_0/D ypass vdd vdd pmos_3p3 w=1.485u l=0.6u
X1 vdd ypass nmos_5p0431058998322_64x8m81_0/D vdd pmos_3p3 w=1.485u l=0.6u
X2 a_447_11191# pcb a_222_11191# vdd pmos_3p3 w=3.41u l=0.6u
X3 a_222_11191# pcb a_n4_11191# vdd pmos_3p3 w=3.41u l=0.6u
X4 a_447_10416# pcb a_222_10416# vdd pmos_3p3 w=3.41u l=0.6u
X5 a_222_10416# pcb a_n4_10416# vdd pmos_3p3 w=3.41u l=0.6u
.ends

.subckt ypass_gate_64x8m81 d pcb b bb ypass m3_n1_4331# m3_n1_1708# db m3_n1_1160#
+ m3_n1_2030# vdd m3_n1_3366# m3_n1_2352# m3_n1_3688# m3_n1_4009# vss m3_n1_2674#
Xpmos_5p0431058998321_64x8m81_0 vdd b pcb bb pmos_5p0431058998321_64x8m81
Xpmos_5p0431058998321_64x8m81_1 vdd db nmos_5p0431058998322_64x8m81_0/D bb pmos_5p0431058998321_64x8m81
Xnmos_1p2$$47119404_64x8m81_0 d b ypass vss nmos_1p2$$47119404_64x8m81
Xnmos_1p2$$47119404_64x8m81_1 db bb ypass vss nmos_1p2$$47119404_64x8m81
Xpmos_1p2$$46889004_64x8m81_0 d vdd b nmos_5p0431058998322_64x8m81_0/D pmos_1p2$$46889004_64x8m81
Xnmos_5p0431058998322_64x8m81_0 nmos_5p0431058998322_64x8m81_0/D ypass vss ypass vss
+ nmos_5p0431058998322_64x8m81
X0 nmos_5p0431058998322_64x8m81_0/D ypass vdd vdd pmos_3p3 w=1.485u l=0.6u
X1 vdd pcb bb vdd pmos_3p3 w=3.41u l=0.6u
X2 bb pcb vdd vdd pmos_3p3 w=3.41u l=0.6u
X3 vdd pcb b vdd pmos_3p3 w=3.41u l=0.6u
X4 vdd ypass nmos_5p0431058998322_64x8m81_0/D vdd pmos_3p3 w=1.485u l=0.6u
X5 b pcb vdd vdd pmos_3p3 w=3.41u l=0.6u
.ends

.subckt mux821_64x8m81 a_656_7735# ypass_gate_a_64x8m81_0/a_222_11191# ypass_gate_64x8m81_0/d
+ ypass_gate_64x8m81_4/b ypass_gate_64x8m81_6/m3_n1_1708# ypass_gate_64x8m81_2/d ypass_gate_a_64x8m81_0/a_447_11191#
+ ypass_gate_64x8m81_6/m3_n1_2030# ypass_gate_64x8m81_4/d ypass_gate_64x8m81_6/db
+ ypass_gate_64x8m81_4/db ypass_gate_64x8m81_6/m3_n1_3366# ypass_gate_64x8m81_6/d
+ ypass_gate_64x8m81_6/m3_n1_2352# ypass_gate_64x8m81_0/ypass ypass_gate_64x8m81_1/ypass
+ ypass_gate_64x8m81_2/ypass ypass_gate_64x8m81_6/m3_n1_3688# ypass_gate_a_64x8m81_0/d
+ ypass_gate_64x8m81_6/m3_n1_4009# ypass_gate_a_64x8m81_0/ypass ypass_gate_64x8m81_3/ypass
+ ypass_gate_a_64x8m81_0/a_222_10416# ypass_gate_64x8m81_6/m3_n1_2674# ypass_gate_a_64x8m81_0/b
+ ypass_gate_64x8m81_4/ypass ypass_gate_64x8m81_5/ypass ypass_gate_64x8m81_6/ypass
+ ypass_gate_64x8m81_1/d ypass_gate_64x8m81_5/db a_4992_424# ypass_gate_a_64x8m81_0/a_447_10416#
+ ypass_gate_64x8m81_3/d ypass_gate_a_64x8m81_0/a_n80_n10# ypass_gate_64x8m81_6/vdd
+ ypass_gate_a_64x8m81_0/db ypass_gate_64x8m81_5/d ypass_gate_64x8m81_6/vss ypass_gate_64x8m81_6/pcb
+ ypass_gate_64x8m81_6/m3_n1_4331#
Xypass_gate_a_64x8m81_0 ypass_gate_a_64x8m81_0/d ypass_gate_64x8m81_6/pcb ypass_gate_64x8m81_6/vss
+ ypass_gate_a_64x8m81_0/b ypass_gate_a_64x8m81_0/bb ypass_gate_a_64x8m81_0/db ypass_gate_a_64x8m81_0/ypass
+ ypass_gate_a_64x8m81_0/a_222_11191# ypass_gate_64x8m81_6/vdd ypass_gate_64x8m81_6/m3_n1_4331#
+ ypass_gate_a_64x8m81_0/a_447_11191# ypass_gate_a_64x8m81_0/a_n80_n10# ypass_gate_a_64x8m81_0/a_222_10416#
+ ypass_gate_64x8m81_6/m3_n1_1708# ypass_gate_64x8m81_6/vdd ypass_gate_64x8m81_6/vdd
+ ypass_gate_64x8m81_6/m3_n1_2030# ypass_gate_64x8m81_6/vdd ypass_gate_64x8m81_1/db
+ ypass_gate_64x8m81_6/m3_n1_3366# ypass_gate_a_64x8m81_0/a_447_10416# ypass_gate_64x8m81_6/m3_n1_2352#
+ ypass_gate_64x8m81_6/m3_n1_3688# ypass_gate_64x8m81_6/m3_n1_4009# ypass_gate_64x8m81_6/m3_n1_2674#
+ ypass_gate_a_64x8m81
Xypass_gate_64x8m81_1 ypass_gate_64x8m81_1/d ypass_gate_64x8m81_6/pcb ypass_gate_64x8m81_1/b
+ ypass_gate_64x8m81_1/bb ypass_gate_64x8m81_1/ypass ypass_gate_64x8m81_6/m3_n1_4331#
+ ypass_gate_64x8m81_6/m3_n1_1708# ypass_gate_64x8m81_1/db ypass_gate_64x8m81_6/vdd
+ ypass_gate_64x8m81_6/m3_n1_2030# ypass_gate_64x8m81_6/vdd ypass_gate_64x8m81_6/m3_n1_3366#
+ ypass_gate_64x8m81_6/m3_n1_2352# ypass_gate_64x8m81_6/m3_n1_3688# ypass_gate_64x8m81_6/m3_n1_4009#
+ ypass_gate_64x8m81_6/vss ypass_gate_64x8m81_6/m3_n1_2674# ypass_gate_64x8m81
Xypass_gate_64x8m81_0 ypass_gate_64x8m81_0/d ypass_gate_64x8m81_6/pcb ypass_gate_64x8m81_0/b
+ ypass_gate_64x8m81_0/bb ypass_gate_64x8m81_0/ypass ypass_gate_64x8m81_6/m3_n1_4331#
+ ypass_gate_64x8m81_6/m3_n1_1708# ypass_gate_64x8m81_4/db ypass_gate_64x8m81_6/vdd
+ ypass_gate_64x8m81_6/m3_n1_2030# ypass_gate_64x8m81_6/vdd ypass_gate_64x8m81_6/m3_n1_3366#
+ ypass_gate_64x8m81_6/m3_n1_2352# ypass_gate_64x8m81_6/m3_n1_3688# ypass_gate_64x8m81_6/m3_n1_4009#
+ ypass_gate_64x8m81_6/vss ypass_gate_64x8m81_6/m3_n1_2674# ypass_gate_64x8m81
Xypass_gate_64x8m81_2 ypass_gate_64x8m81_2/d ypass_gate_64x8m81_6/pcb ypass_gate_64x8m81_2/b
+ ypass_gate_64x8m81_2/bb ypass_gate_64x8m81_2/ypass ypass_gate_64x8m81_6/m3_n1_4331#
+ ypass_gate_64x8m81_6/m3_n1_1708# ypass_gate_64x8m81_5/db ypass_gate_64x8m81_6/vdd
+ ypass_gate_64x8m81_6/m3_n1_2030# ypass_gate_64x8m81_6/vdd ypass_gate_64x8m81_6/m3_n1_3366#
+ ypass_gate_64x8m81_6/m3_n1_2352# ypass_gate_64x8m81_6/m3_n1_3688# ypass_gate_64x8m81_6/m3_n1_4009#
+ ypass_gate_64x8m81_6/vss ypass_gate_64x8m81_6/m3_n1_2674# ypass_gate_64x8m81
Xypass_gate_64x8m81_3 ypass_gate_64x8m81_3/d ypass_gate_64x8m81_6/pcb ypass_gate_64x8m81_3/b
+ ypass_gate_64x8m81_3/bb ypass_gate_64x8m81_3/ypass ypass_gate_64x8m81_6/m3_n1_4331#
+ ypass_gate_64x8m81_6/m3_n1_1708# ypass_gate_64x8m81_6/db ypass_gate_64x8m81_6/vdd
+ ypass_gate_64x8m81_6/m3_n1_2030# ypass_gate_64x8m81_6/vdd ypass_gate_64x8m81_6/m3_n1_3366#
+ ypass_gate_64x8m81_6/m3_n1_2352# ypass_gate_64x8m81_6/m3_n1_3688# ypass_gate_64x8m81_6/m3_n1_4009#
+ ypass_gate_64x8m81_6/vss ypass_gate_64x8m81_6/m3_n1_2674# ypass_gate_64x8m81
Xypass_gate_64x8m81_4 ypass_gate_64x8m81_4/d ypass_gate_64x8m81_6/pcb ypass_gate_64x8m81_4/b
+ ypass_gate_64x8m81_4/bb ypass_gate_64x8m81_4/ypass ypass_gate_64x8m81_6/m3_n1_4331#
+ ypass_gate_64x8m81_6/m3_n1_1708# ypass_gate_64x8m81_4/db ypass_gate_64x8m81_6/vdd
+ ypass_gate_64x8m81_6/m3_n1_2030# ypass_gate_64x8m81_6/vdd ypass_gate_64x8m81_6/m3_n1_3366#
+ ypass_gate_64x8m81_6/m3_n1_2352# ypass_gate_64x8m81_6/m3_n1_3688# ypass_gate_64x8m81_6/m3_n1_4009#
+ ypass_gate_64x8m81_6/vss ypass_gate_64x8m81_6/m3_n1_2674# ypass_gate_64x8m81
Xypass_gate_64x8m81_5 ypass_gate_64x8m81_5/d ypass_gate_64x8m81_6/pcb ypass_gate_64x8m81_5/b
+ ypass_gate_64x8m81_5/bb ypass_gate_64x8m81_5/ypass ypass_gate_64x8m81_6/m3_n1_4331#
+ ypass_gate_64x8m81_6/m3_n1_1708# ypass_gate_64x8m81_5/db ypass_gate_64x8m81_6/vdd
+ ypass_gate_64x8m81_6/m3_n1_2030# ypass_gate_64x8m81_6/vdd ypass_gate_64x8m81_6/m3_n1_3366#
+ ypass_gate_64x8m81_6/m3_n1_2352# ypass_gate_64x8m81_6/m3_n1_3688# ypass_gate_64x8m81_6/m3_n1_4009#
+ ypass_gate_64x8m81_6/vss ypass_gate_64x8m81_6/m3_n1_2674# ypass_gate_64x8m81
Xypass_gate_64x8m81_6 ypass_gate_64x8m81_6/d ypass_gate_64x8m81_6/pcb ypass_gate_64x8m81_6/b
+ ypass_gate_64x8m81_6/bb ypass_gate_64x8m81_6/ypass ypass_gate_64x8m81_6/m3_n1_4331#
+ ypass_gate_64x8m81_6/m3_n1_1708# ypass_gate_64x8m81_6/db ypass_gate_64x8m81_6/vdd
+ ypass_gate_64x8m81_6/m3_n1_2030# ypass_gate_64x8m81_6/vdd ypass_gate_64x8m81_6/m3_n1_3366#
+ ypass_gate_64x8m81_6/m3_n1_2352# ypass_gate_64x8m81_6/m3_n1_3688# ypass_gate_64x8m81_6/m3_n1_4009#
+ ypass_gate_64x8m81_6/vss ypass_gate_64x8m81_6/m3_n1_2674# ypass_gate_64x8m81
.ends

.subckt saout_R_m2_64x8m81 pcb datain WEN ypass[1] ypass[2] ypass[3] ypass[4] ypass[5]
+ ypass[6] ypass[7] men ypass[0] GWEN b[0] q bb[1] sa_64x8m81_0/wep outbuf_oe_64x8m81_0/a_4913_n316#
+ GWE bb[2] b[3] bb[5] mux821_64x8m81_0/ypass_gate_a_64x8m81_0/ypass bb[0] sacntl_2_64x8m81_0/a_4560_1922#
+ mux821_64x8m81_0/a_656_7735# b[7] wen_wm1_64x8m81_0/GWEN a_5189_27169# a_5414_27169#
+ b[2] b[6] bb[3] a_5189_27944# a_5414_27944# b[5] b[1] bb[4] din_64x8m81_0/men b[4]
+ mux821_64x8m81_0/ypass_gate_64x8m81_3/ypass bb[6] mux821_64x8m81_0/ypass_gate_64x8m81_2/ypass
+ mux821_64x8m81_0/ypass_gate_64x8m81_6/ypass wen_wm1_64x8m81_0/wen mux821_64x8m81_0/ypass_gate_64x8m81_4/ypass
+ wen_wm1_64x8m81_0/vdd bb[7] mux821_64x8m81_0/ypass_gate_64x8m81_1/ypass sa_64x8m81_0/pcb
+ sacntl_2_64x8m81_0/a_4718_983# mux821_64x8m81_0/ypass_gate_64x8m81_4/b mux821_64x8m81_0/ypass_gate_64x8m81_5/ypass
+ mux821_64x8m81_0/ypass_gate_64x8m81_0/ypass vss mux821_64x8m81_0/ypass_gate_64x8m81_6/vdd
+ sacntl_2_64x8m81_0/vdd vdd
Xsa_64x8m81_0 sa_64x8m81_0/wep sa_64x8m81_0/se sa_64x8m81_0/pcb sa_64x8m81_0/qp vdd
+ vss sa_64x8m81
Xwen_wm1_64x8m81_0 sa_64x8m81_0/wep wen_wm1_64x8m81_0/wen wen_wm1_64x8m81_0/GWEN vss
+ din_64x8m81_0/men wen_wm1_64x8m81_0/vdd wen_wm1_64x8m81
Xsacntl_2_64x8m81_0 sa_64x8m81_0/pcb sa_64x8m81_0/se din_64x8m81_0/men sacntl_2_64x8m81_0/pmos_1p2$$46282796_64x8m81_0/pmos_5p04310589983223_64x8m81_0/D
+ sacntl_2_64x8m81_0/a_4718_983# vss sacntl_2_64x8m81_0/pmos_5p04310589983226_64x8m81_2/S
+ sacntl_2_64x8m81_0/pmos_5p04310589983226_64x8m81_1/S sacntl_2_64x8m81_0/a_4560_1922#
+ sacntl_2_64x8m81_0/pmos_5p04310589983226_64x8m81_2/S sacntl_2_64x8m81_0/vdd vss
+ sacntl_2_64x8m81
Xoutbuf_oe_64x8m81_0 sa_64x8m81_0/se q GWE sa_64x8m81_0/qp sa_64x8m81_0/qp outbuf_oe_64x8m81_0/a_4913_n316#
+ vdd vss outbuf_oe_64x8m81
Xdin_64x8m81_0 datain sa_64x8m81_0/wep din_64x8m81_0/men vdd vdd vdd sa_64x8m81_0/pcb
+ vdd vss din_64x8m81
Xmux821_64x8m81_0 mux821_64x8m81_0/a_656_7735# a_5189_27944# vdd mux821_64x8m81_0/ypass_gate_64x8m81_4/b
+ mux821_64x8m81_0/ypass_gate_64x8m81_3/ypass vdd a_5414_27944# mux821_64x8m81_0/ypass_gate_64x8m81_6/ypass
+ vdd vdd vdd mux821_64x8m81_0/ypass_gate_64x8m81_0/ypass vdd mux821_64x8m81_0/ypass_gate_64x8m81_2/ypass
+ mux821_64x8m81_0/ypass_gate_64x8m81_0/ypass mux821_64x8m81_0/ypass_gate_64x8m81_1/ypass
+ mux821_64x8m81_0/ypass_gate_64x8m81_2/ypass mux821_64x8m81_0/ypass_gate_64x8m81_4/ypass
+ vdd mux821_64x8m81_0/ypass_gate_64x8m81_1/ypass mux821_64x8m81_0/ypass_gate_a_64x8m81_0/ypass
+ mux821_64x8m81_0/ypass_gate_64x8m81_3/ypass a_5189_27169# mux821_64x8m81_0/ypass_gate_64x8m81_5/ypass
+ mux821_64x8m81_0/ypass_gate_a_64x8m81_0/b mux821_64x8m81_0/ypass_gate_64x8m81_4/ypass
+ mux821_64x8m81_0/ypass_gate_64x8m81_5/ypass mux821_64x8m81_0/ypass_gate_64x8m81_6/ypass
+ vdd vdd mux821_64x8m81_0/a_4992_424# a_5414_27169# vdd mux821_64x8m81_0/ypass_gate_a_64x8m81_0/a_n80_n10#
+ mux821_64x8m81_0/ypass_gate_64x8m81_6/vdd vdd vdd vss sa_64x8m81_0/pcb mux821_64x8m81_0/ypass_gate_a_64x8m81_0/ypass
+ mux821_64x8m81
.ends

.subckt x018SRAM_cell1_64x8m81 a_n36_52# a_444_n42# a_246_342# a_246_712# m3_n36_330#
+ a_36_n42# w_n68_622# VSUBS
X0 a_126_298# a_n36_52# a_444_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X1 a_36_206# a_n36_52# a_36_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X2 a_246_712# a_126_298# a_36_206# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X3 a_126_298# a_36_206# a_246_712# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X4 a_246_342# a_126_298# a_36_206# VSUBS nmos_6p0 w=0.95u l=0.6u
X5 a_126_298# a_36_206# a_246_342# VSUBS nmos_6p0 w=0.95u l=0.6u
.ends

.subckt x018SRAM_cell1_2x_64x8m81 018SRAM_cell1_64x8m81_1/m3_n36_330# 018SRAM_cell1_64x8m81_0/m3_n36_330#
+ 018SRAM_cell1_64x8m81_0/a_246_342# 018SRAM_cell1_64x8m81_0/a_246_712# 018SRAM_cell1_64x8m81_1/a_444_n42#
+ 018SRAM_cell1_64x8m81_1/a_246_342# 018SRAM_cell1_64x8m81_1/a_246_712# 018SRAM_cell1_64x8m81_1/a_36_n42#
+ 018SRAM_cell1_64x8m81_0/a_n36_52# 018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_64x8m81_0/w_n68_622#
+ 018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS
X018SRAM_cell1_64x8m81_0 018SRAM_cell1_64x8m81_0/a_n36_52# 018SRAM_cell1_64x8m81_1/a_444_n42#
+ 018SRAM_cell1_64x8m81_0/a_246_342# 018SRAM_cell1_64x8m81_0/a_246_712# 018SRAM_cell1_64x8m81_0/m3_n36_330#
+ 018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_64x8m81
X018SRAM_cell1_64x8m81_1 018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_64x8m81_1/a_444_n42#
+ 018SRAM_cell1_64x8m81_1/a_246_342# 018SRAM_cell1_64x8m81_1/a_246_712# 018SRAM_cell1_64x8m81_1/m3_n36_330#
+ 018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_64x8m81
.ends

.subckt col_64a_64x8m81 WL[0] WL[6] WL[4] WL[3] WL[7] WL[1] 018SRAM_cell1_2x_64x8m81_5/018SRAM_cell1_64x8m81_1/a_444_n42#
+ b[5] 018SRAM_cell1_2x_64x8m81_37/018SRAM_cell1_64x8m81_1/a_444_n42# b[1] 018SRAM_cell1_2x_64x8m81_89/018SRAM_cell1_64x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_64x8m81_91/018SRAM_cell1_64x8m81_1/a_444_n42# b[7] 018SRAM_cell1_2x_64x8m81_90/018SRAM_cell1_64x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_64x8m81_4/018SRAM_cell1_64x8m81_1/a_444_n42# WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_64x8m81_98/018SRAM_cell1_64x8m81_1/a_444_n42# b[3] 018SRAM_cell1_2x_64x8m81_80/018SRAM_cell1_64x8m81_1/a_444_n42#
+ bb[4] b[6] 018SRAM_cell1_2x_64x8m81_76/018SRAM_cell1_64x8m81_1/a_444_n42# b[4] 018SRAM_cell1_2x_64x8m81_94/018SRAM_cell1_64x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_64x8m81_1/018SRAM_cell1_64x8m81_1/a_444_n42# WL[2] 018SRAM_cell1_2x_64x8m81_35/018SRAM_cell1_64x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_444_n42# BL bb[7] BL1B 018SRAM_cell1_2x_64x8m81_39/018SRAM_cell1_64x8m81_1/a_444_n42#
+ VSS b[0] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
X018SRAM_cell1_2x_64x8m81_1 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_1/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[0] WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_2 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[0]
+ WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_3 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# b[0] WL[0]
+ WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_4 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_4/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ b[3] WL[0] WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_5 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_5/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[0] WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_6 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[0]
+ WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_7 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ bb[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# b[4] WL[0]
+ WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_8 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[0]
+ WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_9 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ b[5] WL[0] WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_90 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_90/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[2] WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_91 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_91/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[4] WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_80 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_80/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[4] WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_92 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_1/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[4] WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_70 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_5/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[4] WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_81 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_89/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[4] WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_120 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_35/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[4] WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_60 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[6]
+ WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_82 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[2]
+ WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_93 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[4]
+ WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_71 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[4]
+ WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_110 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# b[0] WL[2]
+ WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_121 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[4]
+ WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_61 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[6]
+ WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_50 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_98/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ b[1] WL[6] WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_94 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_94/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[4] WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_83 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_94/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[2] WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_72 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[4]
+ WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_122 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[4]
+ WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_100 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[2]
+ WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_111 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[2]
+ WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_51 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_1/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[6] WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_62 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# b[6] WL[6]
+ WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_40 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_89/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[6] WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_95 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[4]
+ WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_73 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[2]
+ WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_84 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[2]
+ WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_101 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_37/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[2] WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_112 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_4/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ b[3] WL[2] WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_123 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_37/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[4] WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_63 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[6]
+ WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_52 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ b[5] WL[6] WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_41 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_80/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[6] WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_74 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_91/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[2] WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_30 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[0]
+ WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_96 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ bb[7] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# b[7] WL[2]
+ WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_85 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_5/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[2] WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_102 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[2]
+ WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_113 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ bb[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# b[4] WL[2]
+ WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_124 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[4]
+ WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_20 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_76/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[0] WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_53 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_5/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[6] WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_42 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_91/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[6] WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_64 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[4]
+ WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_97 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# b[0] WL[4]
+ WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_75 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[2]
+ WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_31 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_80/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[0] WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_86 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[2]
+ WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_125 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ b[5] WL[4] WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_103 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_35/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[2] WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_114 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ b[5] WL[2] WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_54 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_94/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[6] WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_43 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[6]
+ WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_32 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[6]
+ WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_65 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[4]
+ WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_98 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_98/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ b[1] WL[4] WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_21 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_35/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[0] WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_76 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_76/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[2] WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_10 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_98/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ b[1] WL[0] WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_87 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_1/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[2] WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_104 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[2]
+ WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_115 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# b[6] WL[2]
+ WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_126 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[4] WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_55 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ bb[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# b[4] WL[6]
+ WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_44 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[6]
+ WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_33 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[6]
+ WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_66 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[4]
+ WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_99 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[2] WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_22 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[0] WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_77 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[2]
+ WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_11 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_90/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[0] WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_88 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[2]
+ WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_116 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ bb[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# b[4] WL[4]
+ WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_127 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# b[6] WL[4]
+ WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_105 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[2]
+ WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_56 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[6]
+ WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_45 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[6]
+ WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_34 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[6] WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_23 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[0]
+ WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_78 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_80/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[2] WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_89 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_89/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[2] WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_12 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_94/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[0] WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_67 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_76/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[4] WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_106 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_4/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ b[3] WL[4] WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_117 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_39/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[4] WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_57 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_4/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ b[3] WL[6] WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_46 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_76/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[6] WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_35 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_35/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[6] WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_24 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[0]
+ WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_79 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[2]
+ WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_13 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# b[6] WL[0]
+ WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_68 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[4]
+ WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_107 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_39/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[2] WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_118 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[4]
+ WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_58 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ bb[7] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# b[7] WL[6]
+ WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_36 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[6]
+ WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_47 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[6]
+ WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_69 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_90/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[4] WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_25 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[0]
+ WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_14 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ bb[7] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# b[7] WL[0]
+ WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_108 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ bb[7] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# b[7] WL[4]
+ WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_119 WL[5] WL[4] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[4]
+ WL[5] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_48 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[6]
+ WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_59 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# b[0] WL[6]
+ WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_37 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_37/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[6] WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_26 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_89/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[0] WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_15 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[0]
+ WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_109 WL[3] WL[2] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_98/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ b[1] WL[2] WL[3] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_49 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_90/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[6] WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_38 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[6]
+ WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_16 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_37/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[0] WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_27 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[0]
+ WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_39 WL[7] WL[6] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_39/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[6] WL[7] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_28 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[0]
+ WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_17 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[0]
+ WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_18 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_91/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[0] WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_29 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[0]
+ WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_19 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_39/018SRAM_cell1_64x8m81_1/a_444_n42# VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL WL[0] WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_0 WL[1] WL[0] VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ BL1B VSS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# BL WL[0]
+ WL[1] 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSS x018SRAM_cell1_2x_64x8m81
.ends

.subckt saout_m2_64x8m81 pcb datain WEN ypass[1] ypass[2] ypass[3] ypass[4] ypass[5]
+ ypass[6] ypass[7] men ypass[0] GWEN bb[5] bb[6] b[0] q a_5189_27176# a_5414_27176#
+ sa_64x8m81_0/wep a_5189_27951# a_5414_27951# outbuf_oe_64x8m81_0/a_4913_n316# GWE
+ mux821_64x8m81_0/a_4992_424# b[4] bb[2] bb[7] sacntl_2_64x8m81_0/a_4560_1922# mux821_64x8m81_0/a_656_7735#
+ wen_wm1_64x8m81_0/GWEN mux821_64x8m81_0/ypass_gate_64x8m81_3/ypass b[7] b[5] b[1]
+ bb[4] b[2] b[6] bb[3] b[3] mux821_64x8m81_0/ypass_gate_a_64x8m81_0/a_n80_n10# mux821_64x8m81_0/ypass_gate_a_64x8m81_0/ypass
+ bb[1] mux821_64x8m81_0/ypass_gate_64x8m81_4/ypass mux821_64x8m81_0/ypass_gate_64x8m81_1/ypass
+ wen_wm1_64x8m81_0/vdd bb[0] sa_64x8m81_0/pcb sacntl_2_64x8m81_0/a_4718_983# din_64x8m81_0/men
+ mux821_64x8m81_0/ypass_gate_64x8m81_2/ypass sacntl_2_64x8m81_0/vdd mux821_64x8m81_0/ypass_gate_64x8m81_0/ypass
+ mux821_64x8m81_0/ypass_gate_64x8m81_5/ypass mux821_64x8m81_0/ypass_gate_a_64x8m81_0/b
+ mux821_64x8m81_0/ypass_gate_64x8m81_6/ypass vss mux821_64x8m81_0/ypass_gate_64x8m81_6/vdd
+ vdd
Xsa_64x8m81_0 sa_64x8m81_0/wep sa_64x8m81_0/se sa_64x8m81_0/pcb sa_64x8m81_0/qp vdd
+ vss sa_64x8m81
Xwen_wm1_64x8m81_0 sa_64x8m81_0/wep wen_wm1_64x8m81_0/wen wen_wm1_64x8m81_0/GWEN vss
+ din_64x8m81_0/men wen_wm1_64x8m81_0/vdd wen_wm1_64x8m81
Xsacntl_2_64x8m81_0 sa_64x8m81_0/pcb sa_64x8m81_0/se din_64x8m81_0/men sacntl_2_64x8m81_0/pmos_1p2$$46282796_64x8m81_0/pmos_5p04310589983223_64x8m81_0/D
+ sacntl_2_64x8m81_0/a_4718_983# vss sacntl_2_64x8m81_0/pmos_5p04310589983226_64x8m81_2/S
+ sacntl_2_64x8m81_0/pmos_5p04310589983226_64x8m81_1/S sacntl_2_64x8m81_0/a_4560_1922#
+ sacntl_2_64x8m81_0/pmos_5p04310589983226_64x8m81_2/S sacntl_2_64x8m81_0/vdd vss
+ sacntl_2_64x8m81
Xoutbuf_oe_64x8m81_0 sa_64x8m81_0/se q GWE sa_64x8m81_0/qp sa_64x8m81_0/qp outbuf_oe_64x8m81_0/a_4913_n316#
+ vdd vss outbuf_oe_64x8m81
Xdin_64x8m81_0 datain sa_64x8m81_0/wep din_64x8m81_0/men vdd vdd vdd sa_64x8m81_0/pcb
+ vdd vss din_64x8m81
Xmux821_64x8m81_0 mux821_64x8m81_0/a_656_7735# a_5189_27951# vdd mux821_64x8m81_0/ypass_gate_64x8m81_4/b
+ mux821_64x8m81_0/ypass_gate_a_64x8m81_0/ypass vdd a_5414_27951# mux821_64x8m81_0/ypass_gate_64x8m81_1/ypass
+ vdd vdd vdd mux821_64x8m81_0/ypass_gate_64x8m81_5/ypass vdd mux821_64x8m81_0/ypass_gate_64x8m81_4/ypass
+ mux821_64x8m81_0/ypass_gate_64x8m81_0/ypass mux821_64x8m81_0/ypass_gate_64x8m81_1/ypass
+ mux821_64x8m81_0/ypass_gate_64x8m81_2/ypass mux821_64x8m81_0/ypass_gate_64x8m81_2/ypass
+ vdd mux821_64x8m81_0/ypass_gate_64x8m81_6/ypass mux821_64x8m81_0/ypass_gate_a_64x8m81_0/ypass
+ mux821_64x8m81_0/ypass_gate_64x8m81_3/ypass a_5189_27176# mux821_64x8m81_0/ypass_gate_64x8m81_0/ypass
+ mux821_64x8m81_0/ypass_gate_a_64x8m81_0/b mux821_64x8m81_0/ypass_gate_64x8m81_4/ypass
+ mux821_64x8m81_0/ypass_gate_64x8m81_5/ypass mux821_64x8m81_0/ypass_gate_64x8m81_6/ypass
+ vdd vdd mux821_64x8m81_0/a_4992_424# a_5414_27176# vdd mux821_64x8m81_0/ypass_gate_a_64x8m81_0/a_n80_n10#
+ mux821_64x8m81_0/ypass_gate_64x8m81_6/vdd vdd vdd vss sa_64x8m81_0/pcb mux821_64x8m81_0/ypass_gate_64x8m81_3/ypass
+ mux821_64x8m81
.ends

.subckt x018SRAM_cell1_dummy_R_64x8m81 a_n36_52# a_444_n42# a_246_342# a_126_298#
+ m3_n36_330# a_36_n42# w_n68_622# VSUBS
X0 a_444_206# a_n36_52# a_444_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X1 a_36_206# a_n36_52# a_36_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X2 a_126_298# a_126_298# a_36_206# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X3 a_444_206# a_246_342# a_126_298# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X4 a_246_342# a_126_298# a_36_206# VSUBS nmos_6p0 w=0.95u l=0.6u
X5 a_444_206# a_246_342# a_246_342# VSUBS nmos_6p0 w=0.95u l=0.6u
.ends

.subckt ypass_gate_64x8m81_0 d pcb vss bb db ypass vdd pmos_5p0431058998321_64x8m81_2/D
+ m3_n1_4331# m3_n1_1708# m3_n1_1160# m3_n1_2030# m3_n1_3366# b m3_n1_2352# m3_n1_3688#
+ m3_n1_4009# m3_n1_2674# a_66_539#
Xnmos_5p0431058998320_64x8m81_0 pmos_5p0431058998321_64x8m81_2/D a_66_539# bb vss
+ nmos_5p0431058998320_64x8m81
Xnmos_5p0431058998320_64x8m81_1 d a_66_539# b vss nmos_5p0431058998320_64x8m81
Xpmos_5p0431058998321_64x8m81_0 vdd d nmos_5p0431058998322_64x8m81_0/D b pmos_5p0431058998321_64x8m81
Xpmos_5p0431058998321_64x8m81_1 vdd b pcb bb pmos_5p0431058998321_64x8m81
Xpmos_5p0431058998321_64x8m81_2 vdd pmos_5p0431058998321_64x8m81_2/D nmos_5p0431058998322_64x8m81_0/D
+ bb pmos_5p0431058998321_64x8m81
Xnmos_5p0431058998322_64x8m81_0 nmos_5p0431058998322_64x8m81_0/D a_66_539# vss a_66_539#
+ vss nmos_5p0431058998322_64x8m81
X0 nmos_5p0431058998322_64x8m81_0/D a_66_539# vdd vdd pmos_3p3 w=1.485u l=0.6u
X1 vdd pcb bb vdd pmos_3p3 w=3.41u l=0.6u
X2 bb pcb vdd vdd pmos_3p3 w=3.41u l=0.6u
X3 vdd pcb b vdd pmos_3p3 w=3.41u l=0.6u
X4 vdd a_66_539# nmos_5p0431058998322_64x8m81_0/D vdd pmos_3p3 w=1.485u l=0.6u
X5 b pcb vdd vdd pmos_3p3 w=3.41u l=0.6u
.ends

.subckt x018SRAM_cell1_dummy_64x8m81 a_n36_52# m2_90_n50# a_246_342# m2_390_n50# a_246_712#
+ m3_n36_330# w_n68_622# VSUBS
X0 a_126_298# a_n36_52# a_444_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X1 a_36_206# a_n36_52# a_36_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X2 a_246_712# a_126_298# a_36_206# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X3 a_126_298# a_36_206# a_246_712# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X4 a_246_342# a_126_298# a_36_206# VSUBS nmos_6p0 w=0.95u l=0.6u
X5 a_126_298# a_36_206# a_246_342# VSUBS nmos_6p0 w=0.95u l=0.6u
.ends

.subckt pmos_5p04310589983254_64x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=3.51u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=3.51u l=0.6u
.ends

.subckt new_dummyrow_unit_64x8m81 018SRAM_cell1_dummy_64x8m81_12/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_4/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_13/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_5/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_14/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_6/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_15/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_7/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_8/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_9/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_0/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_2/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_1/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_3/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_4/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_5/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_6/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_7/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_8/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_10/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_9/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_0/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_11/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_13/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_12/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_14/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_1/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_15/m2_390_n50#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_10/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_2/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_11/m2_90_n50# VSUBS 018SRAM_cell1_dummy_64x8m81_3/m2_90_n50#
+ 018SRAM_strap1_64x8m81_1/w_n68_622#
X018SRAM_cell1_dummy_64x8m81_10 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_10/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_10/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_11 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_11/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_11/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_12 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_12/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_12/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_13 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_13/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_13/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_14 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_14/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_14/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_15 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_15/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_15/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_0 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_0/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_0/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_1 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_1/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_1/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_2 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_2/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_2/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_3 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_3/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_3/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_5 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_5/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_5/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_4 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_4/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_4/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_6 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_6/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_6/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_7 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_7/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_7/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_8 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_8/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_8/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_9 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_9/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_9/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
.ends

.subckt nmos_5p04310589983253_64x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=8.5u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=8.5u l=0.6u
.ends

.subckt pmos_5p04310589983255_64x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=10.64u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=10.64u l=0.6u
.ends

.subckt nmos_5p04310589983256_64x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=1.38u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=1.38u l=0.6u
.ends

.subckt rdummy_64x4_64x8m81 tblhl pcb new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_2/m2_390_n50#
+ m3_22279_n11418# 018SRAM_cell1_dummy_64x8m81_41/m2_90_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_3/m2_390_n50#
+ 018SRAM_cell1_dummy_R_64x8m81_3/a_246_342# 018SRAM_cell1_dummy_64x8m81_12/m2_90_n50#
+ 018SRAM_cell1_dummy_R_64x8m81_0/m3_n36_330# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_4/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_22/m2_90_n50# ypass_gate_64x8m81_0_0/b 018SRAM_cell1_dummy_R_64x8m81_1/m3_n36_330#
+ 018SRAM_cell1_dummy_64x8m81_4/m2_90_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_5/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_32/m2_90_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_6/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_0/m2_90_n50# 018SRAM_cell1_dummy_R_64x8m81_7/a_126_298#
+ 018SRAM_cell1_dummy_64x8m81_42/m2_90_n50# 018SRAM_cell1_dummy_R_64x8m81_3/m3_n36_330#
+ m3_22279_n9439# 018SRAM_cell1_dummy_64x8m81_40/m2_390_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_7/m2_390_n50#
+ m3_22426_n25051# 018SRAM_cell1_dummy_R_64x8m81_4/a_246_342# 018SRAM_cell1_dummy_64x8m81_41/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_13/m2_90_n50# 018SRAM_cell1_dummy_R_64x8m81_4/m3_n36_330#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_8/m2_390_n50# 018SRAM_cell1_2x_64x8m81_1/018SRAM_cell1_64x8m81_1/m3_n36_330#
+ 018SRAM_cell1_dummy_64x8m81_23/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_42/m2_390_n50#
+ 018SRAM_cell1_dummy_R_64x8m81_5/m3_n36_330# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_9/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_5/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_43/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_33/m2_90_n50# 018SRAM_cell1_dummy_R_64x8m81_6/m3_n36_330#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_1/m2_90_n50# 018SRAM_cell1_2x_64x8m81_3/018SRAM_cell1_64x8m81_0/m3_n36_330#
+ 018SRAM_cell1_dummy_64x8m81_43/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_44/m2_390_n50#
+ 018SRAM_cell1_dummy_R_64x8m81_7/m3_n36_330# 018SRAM_cell1_dummy_R_64x8m81_5/a_246_342#
+ 018SRAM_cell1_dummy_64x8m81_45/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_14/m2_90_n50#
+ 018SRAM_cell1_dummy_R_64x8m81_8/m3_n36_330# 018SRAM_cell1_dummy_64x8m81_24/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_46/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_6/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_34/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_47/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_2/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_44/m2_90_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_10/m2_90_n50# 018SRAM_cell1_dummy_R_64x8m81_6/a_246_342#
+ 018SRAM_cell1_dummy_64x8m81_30/m2_390_n50# DWL 018SRAM_cell1_dummy_64x8m81_15/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_25/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_31/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_10/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_7/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_32/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_35/m2_90_n50#
+ a_23395_52# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_3/m2_90_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_11/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_33/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_45/m2_90_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_11/m2_90_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_12/m2_390_n50# 018SRAM_cell1_dummy_R_64x8m81_7/a_246_342#
+ 018SRAM_cell1_dummy_64x8m81_16/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_34/m2_390_n50#
+ m3_22279_n11740# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_13/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_26/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_35/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_14/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_8/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_36/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_36/m2_90_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_15/m2_390_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_4/m2_90_n50#
+ 018SRAM_cell1_dummy_R_64x8m81_5/a_126_298# 018SRAM_cell1_dummy_64x8m81_37/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_46/m2_90_n50# m3_22279_n9760# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_12/m2_90_n50#
+ 018SRAM_cell1_dummy_R_64x8m81_8/a_246_342# 018SRAM_cell1_dummy_64x8m81_17/m2_90_n50#
+ 018SRAM_cell1_2x_64x8m81_3/018SRAM_cell1_64x8m81_1/m3_n36_330# 018SRAM_cell1_dummy_64x8m81_38/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_39/m2_390_n50# 018SRAM_cell1_2x_64x8m81_0/018SRAM_cell1_64x8m81_0/m3_n36_330#
+ 018SRAM_cell1_dummy_64x8m81_20/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_27/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_0/m2_390_n50# 018SRAM_cell1_2x_64x8m81_2/018SRAM_cell1_64x8m81_0/m3_n36_330#
+ 018SRAM_cell1_dummy_64x8m81_9/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_21/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_1/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_37/m2_90_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_5/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_22/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_47/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_2/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_13/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_23/m2_390_n50#
+ 018SRAM_cell1_dummy_R_64x8m81_5/w_n68_622# a_23341_1594# 018SRAM_cell1_dummy_64x8m81_18/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_3/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_24/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_28/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_4/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_25/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_5/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_38/m2_90_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_6/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_26/m2_390_n50# w_22685_n22093# 018SRAM_cell1_dummy_64x8m81_6/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_14/m2_90_n50# m3_22279_n11096#
+ 018SRAM_cell1_dummy_64x8m81_27/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_19/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_7/m2_390_n50# pmos_5p04310589983255_64x8m81_0/S 018SRAM_cell1_dummy_64x8m81_28/m2_390_n50#
+ ypass_gate_64x8m81_0_0/d 018SRAM_cell1_dummy_64x8m81_29/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_8/m2_390_n50#
+ m3_22279_n10082# 018SRAM_cell1_dummy_64x8m81_0/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_29/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_10/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_9/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_39/m2_90_n50# vdd new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_7/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_11/m2_390_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_15/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_12/m2_390_n50# 018SRAM_cell1_dummy_R_64x8m81_0/a_246_342#
+ 018SRAM_cell1_dummy_64x8m81_13/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_1/m2_90_n50#
+ 018SRAM_cell1_2x_64x8m81_0/018SRAM_cell1_64x8m81_1/m3_n36_330# VSS 018SRAM_cell1_dummy_64x8m81_14/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_8/m2_90_n50# 018SRAM_cell1_dummy_R_64x8m81_8/a_126_298#
+ 018SRAM_cell1_dummy_64x8m81_15/m2_390_n50# 018SRAM_cell1_2x_64x8m81_2/018SRAM_cell1_64x8m81_1/m3_n36_330#
+ m3_22279_n10774# 018SRAM_cell1_dummy_R_64x8m81_1/a_246_342# 018SRAM_cell1_2x_64x8m81_1/018SRAM_cell1_64x8m81_0/m3_n36_330#
+ 018SRAM_cell1_dummy_64x8m81_10/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_16/m2_390_n50#
+ 018SRAM_cell1_dummy_R_64x8m81_7/w_n68_622# a_n257_52# 018SRAM_cell1_dummy_64x8m81_20/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_17/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_2/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_18/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_30/m2_90_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_9/m2_90_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_dummy_64x8m81_40/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_19/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_11/m2_90_n50# 018SRAM_cell1_dummy_R_64x8m81_8/w_n68_622#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_0/m2_390_n50# a_n257_1594#
+ 018SRAM_cell1_dummy_64x8m81_21/m2_90_n50# m3_22279_n9117# 018SRAM_cell1_dummy_64x8m81_3/m2_90_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_1/m2_390_n50# vss 018SRAM_cell1_dummy_64x8m81_31/m2_90_n50#
X018SRAM_cell1_2x_64x8m81_1 018SRAM_cell1_2x_64x8m81_1/018SRAM_cell1_64x8m81_1/m3_n36_330#
+ 018SRAM_cell1_2x_64x8m81_1/018SRAM_cell1_64x8m81_0/m3_n36_330# vss 018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_64x8m81_1/a_444_n42# vss 018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_64x8m81_1/a_36_n42#
+ a_n257_1594# a_n257_1594# 018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ vss x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_dummy_R_64x8m81_4 DWL ypass_gate_64x8m81_0_0/bb 018SRAM_cell1_dummy_R_64x8m81_4/a_246_342#
+ 018SRAM_cell1_dummy_R_64x8m81_5/a_126_298# 018SRAM_cell1_dummy_R_64x8m81_4/m3_n36_330#
+ ypass_gate_64x8m81_0_0/b 018SRAM_cell1_dummy_R_64x8m81_5/w_n68_622# vss x018SRAM_cell1_dummy_R_64x8m81
X018SRAM_cell1_2x_64x8m81_2 018SRAM_cell1_2x_64x8m81_2/018SRAM_cell1_64x8m81_1/m3_n36_330#
+ 018SRAM_cell1_2x_64x8m81_2/018SRAM_cell1_64x8m81_0/m3_n36_330# vss 018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_64x8m81_1/a_444_n42# vss 018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_64x8m81_1/a_36_n42#
+ a_n257_1594# a_n257_1594# 018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ vss x018SRAM_cell1_2x_64x8m81
Xypass_gate_64x8m81_0_0 ypass_gate_64x8m81_0_0/d ypass_gate_64x8m81_0_0/pcb vss ypass_gate_64x8m81_0_0/bb
+ ypass_gate_64x8m81_0_0/db ypass_gate_64x8m81_0_0/ypass vdd ypass_gate_64x8m81_0_0/bb
+ m3_22279_n9117# m3_22279_n11740# vdd m3_22279_n11418# m3_22279_n10082# ypass_gate_64x8m81_0_0/b
+ m3_22279_n11096# m3_22279_n9760# m3_22279_n9439# m3_22279_n10774# vdd ypass_gate_64x8m81_0
X018SRAM_cell1_dummy_R_64x8m81_5 a_23341_1594# ypass_gate_64x8m81_0_0/bb 018SRAM_cell1_dummy_R_64x8m81_5/a_246_342#
+ 018SRAM_cell1_dummy_R_64x8m81_5/a_126_298# 018SRAM_cell1_dummy_R_64x8m81_5/m3_n36_330#
+ ypass_gate_64x8m81_0_0/b 018SRAM_cell1_dummy_R_64x8m81_5/w_n68_622# vss x018SRAM_cell1_dummy_R_64x8m81
X018SRAM_cell1_2x_64x8m81_3 018SRAM_cell1_2x_64x8m81_3/018SRAM_cell1_64x8m81_1/m3_n36_330#
+ 018SRAM_cell1_2x_64x8m81_3/018SRAM_cell1_64x8m81_0/m3_n36_330# vss 018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_64x8m81_1/a_444_n42# vss 018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_64x8m81_1/a_36_n42#
+ a_n257_1594# a_n257_1594# 018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ vss x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_dummy_R_64x8m81_6 DWL ypass_gate_64x8m81_0_0/bb 018SRAM_cell1_dummy_R_64x8m81_6/a_246_342#
+ 018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_dummy_R_64x8m81_6/m3_n36_330# ypass_gate_64x8m81_0_0/b
+ 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_R_64x8m81
X018SRAM_cell1_dummy_64x8m81_40 a_n257_52# 018SRAM_cell1_dummy_64x8m81_40/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_40/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_R_64x8m81_7 a_23341_1594# ypass_gate_64x8m81_0_0/bb 018SRAM_cell1_dummy_R_64x8m81_7/a_246_342#
+ 018SRAM_cell1_dummy_R_64x8m81_7/a_126_298# 018SRAM_cell1_dummy_R_64x8m81_7/m3_n36_330#
+ ypass_gate_64x8m81_0_0/b 018SRAM_cell1_dummy_R_64x8m81_7/w_n68_622# vss x018SRAM_cell1_dummy_R_64x8m81
X018SRAM_cell1_dummy_64x8m81_30 DWL 018SRAM_cell1_dummy_64x8m81_30/m2_90_n50# vss
+ 018SRAM_cell1_dummy_64x8m81_30/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622# DWL
+ 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_41 a_n257_52# 018SRAM_cell1_dummy_64x8m81_41/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_41/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_R_64x8m81_8 a_23341_1594# ypass_gate_64x8m81_0_0/bb 018SRAM_cell1_dummy_R_64x8m81_8/a_246_342#
+ 018SRAM_cell1_dummy_R_64x8m81_8/a_126_298# 018SRAM_cell1_dummy_R_64x8m81_8/m3_n36_330#
+ ypass_gate_64x8m81_0_0/b 018SRAM_cell1_dummy_R_64x8m81_8/w_n68_622# vss x018SRAM_cell1_dummy_R_64x8m81
X018SRAM_cell1_dummy_64x8m81_20 DWL 018SRAM_cell1_dummy_64x8m81_20/m2_90_n50# vss
+ 018SRAM_cell1_dummy_64x8m81_20/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622# DWL
+ 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_31 DWL 018SRAM_cell1_dummy_64x8m81_31/m2_90_n50# vss
+ 018SRAM_cell1_dummy_64x8m81_31/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622# DWL
+ 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_42 a_n257_52# 018SRAM_cell1_dummy_64x8m81_42/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_42/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_R_64x8m81_9 a_23395_52# ypass_gate_64x8m81_0_0/bb vss 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# ypass_gate_64x8m81_0_0/b 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_R_64x8m81
X018SRAM_cell1_dummy_64x8m81_43 a_n257_52# 018SRAM_cell1_dummy_64x8m81_43/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_43/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_10 a_n257_52# 018SRAM_cell1_dummy_64x8m81_10/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_10/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_21 DWL 018SRAM_cell1_dummy_64x8m81_21/m2_90_n50# vss
+ 018SRAM_cell1_dummy_64x8m81_21/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622# DWL
+ 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_32 a_n257_52# 018SRAM_cell1_dummy_64x8m81_32/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_32/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
Xpmos_5p04310589983254_64x8m81_0 vdd pmos_5p04310589983254_64x8m81_0/D ypass_gate_64x8m81_0_0/d
+ vdd ypass_gate_64x8m81_0_0/d pmos_5p04310589983254_64x8m81
X018SRAM_cell1_dummy_64x8m81_44 a_n257_52# 018SRAM_cell1_dummy_64x8m81_44/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_44/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_11 a_n257_52# 018SRAM_cell1_dummy_64x8m81_11/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_11/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_22 DWL 018SRAM_cell1_dummy_64x8m81_22/m2_90_n50# vss
+ 018SRAM_cell1_dummy_64x8m81_22/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622# DWL
+ 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_33 a_n257_52# 018SRAM_cell1_dummy_64x8m81_33/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_33/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_45 a_n257_52# 018SRAM_cell1_dummy_64x8m81_45/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_45/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_12 a_n257_52# 018SRAM_cell1_dummy_64x8m81_12/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_12/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_23 DWL 018SRAM_cell1_dummy_64x8m81_23/m2_90_n50# vss
+ 018SRAM_cell1_dummy_64x8m81_23/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622# DWL
+ 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_34 a_n257_52# 018SRAM_cell1_dummy_64x8m81_34/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_34/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_46 a_n257_52# 018SRAM_cell1_dummy_64x8m81_46/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_46/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_13 a_n257_52# 018SRAM_cell1_dummy_64x8m81_13/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_13/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_24 DWL 018SRAM_cell1_dummy_64x8m81_24/m2_90_n50# vss
+ 018SRAM_cell1_dummy_64x8m81_24/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622# DWL
+ 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_35 a_n257_52# 018SRAM_cell1_dummy_64x8m81_35/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_35/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_47 a_n257_52# 018SRAM_cell1_dummy_64x8m81_47/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_47/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_14 a_n257_52# 018SRAM_cell1_dummy_64x8m81_14/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_14/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_25 DWL 018SRAM_cell1_dummy_64x8m81_25/m2_90_n50# vss
+ 018SRAM_cell1_dummy_64x8m81_25/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622# DWL
+ 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_36 a_n257_52# 018SRAM_cell1_dummy_64x8m81_36/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_36/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_15 a_n257_52# 018SRAM_cell1_dummy_64x8m81_15/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_15/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_26 DWL 018SRAM_cell1_dummy_64x8m81_26/m2_90_n50# vss
+ 018SRAM_cell1_dummy_64x8m81_26/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622# DWL
+ 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_37 a_n257_52# 018SRAM_cell1_dummy_64x8m81_37/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_37/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_16 DWL 018SRAM_cell1_dummy_64x8m81_16/m2_90_n50# vss
+ 018SRAM_cell1_dummy_64x8m81_16/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622# DWL
+ 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_27 DWL 018SRAM_cell1_dummy_64x8m81_27/m2_90_n50# vss
+ 018SRAM_cell1_dummy_64x8m81_27/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622# DWL
+ 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_38 a_n257_52# 018SRAM_cell1_dummy_64x8m81_38/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_38/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_0 a_n257_52# 018SRAM_cell1_dummy_64x8m81_0/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_0/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
Xnew_dummyrow_unit_64x8m81_0 new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_12/m2_90_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_4/m2_90_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_13/m2_90_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_5/m2_90_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_14/m2_90_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_6/m2_90_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_15/m2_90_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_7/m2_90_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_8/m2_90_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_9/m2_90_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_0/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_2/m2_390_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_1/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_3/m2_390_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_4/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_5/m2_390_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_6/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_7/m2_390_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_8/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_10/m2_390_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_9/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_0/m2_90_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_11/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_13/m2_390_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_12/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_14/m2_390_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_1/m2_90_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_15/m2_390_n50# DWL new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_10/m2_90_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_2/m2_90_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_11/m2_90_n50#
+ vss new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_3/m2_90_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ new_dummyrow_unit_64x8m81
X018SRAM_cell1_dummy_64x8m81_17 DWL 018SRAM_cell1_dummy_64x8m81_17/m2_90_n50# vss
+ 018SRAM_cell1_dummy_64x8m81_17/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622# DWL
+ 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_28 DWL 018SRAM_cell1_dummy_64x8m81_28/m2_90_n50# vss
+ 018SRAM_cell1_dummy_64x8m81_28/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622# DWL
+ 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_39 a_n257_52# 018SRAM_cell1_dummy_64x8m81_39/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_39/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_1 a_n257_52# 018SRAM_cell1_dummy_64x8m81_1/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_1/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_18 DWL 018SRAM_cell1_dummy_64x8m81_18/m2_90_n50# vss
+ 018SRAM_cell1_dummy_64x8m81_18/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622# DWL
+ 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_29 DWL 018SRAM_cell1_dummy_64x8m81_29/m2_90_n50# vss
+ 018SRAM_cell1_dummy_64x8m81_29/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622# DWL
+ 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_2 a_n257_52# 018SRAM_cell1_dummy_64x8m81_2/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_2/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_3 a_n257_52# 018SRAM_cell1_dummy_64x8m81_3/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_3/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_19 DWL 018SRAM_cell1_dummy_64x8m81_19/m2_90_n50# vss
+ 018SRAM_cell1_dummy_64x8m81_19/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622# DWL
+ 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_64x8m81_0 a_n257_52# 018SRAM_cell1_64x8m81_1/a_444_n42# vss 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ vss x018SRAM_cell1_64x8m81
X018SRAM_cell1_dummy_64x8m81_4 a_n257_52# 018SRAM_cell1_dummy_64x8m81_4/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_4/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_64x8m81_1 a_n257_1594# 018SRAM_cell1_64x8m81_1/a_444_n42# vss 018SRAM_cell1_64x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_64x8m81
X018SRAM_cell1_dummy_64x8m81_5 a_n257_52# 018SRAM_cell1_dummy_64x8m81_5/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_5/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_6 a_n257_52# 018SRAM_cell1_dummy_64x8m81_6/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_6/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_7 a_n257_52# 018SRAM_cell1_dummy_64x8m81_7/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_7/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_8 a_n257_52# 018SRAM_cell1_dummy_64x8m81_8/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_8/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_9 a_n257_52# 018SRAM_cell1_dummy_64x8m81_9/m2_90_n50#
+ vss 018SRAM_cell1_dummy_64x8m81_9/m2_390_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_64x8m81
Xnmos_5p04310589983253_64x8m81_0 tblhl pmos_5p04310589983254_64x8m81_0/D vss pmos_5p04310589983254_64x8m81_0/D
+ vss nmos_5p04310589983253_64x8m81
X018SRAM_cell1_dummy_R_64x8m81_0 a_23341_1594# ypass_gate_64x8m81_0_0/bb 018SRAM_cell1_dummy_R_64x8m81_0/a_246_342#
+ 018SRAM_cell1_dummy_R_64x8m81_7/a_126_298# 018SRAM_cell1_dummy_R_64x8m81_0/m3_n36_330#
+ ypass_gate_64x8m81_0_0/b 018SRAM_cell1_dummy_R_64x8m81_7/w_n68_622# vss x018SRAM_cell1_dummy_R_64x8m81
Xpmos_5p04310589983255_64x8m81_0 w_22685_n22093# tblhl pmos_5p04310589983254_64x8m81_0/D
+ pmos_5p04310589983255_64x8m81_0/S pmos_5p04310589983254_64x8m81_0/D pmos_5p04310589983255_64x8m81
X018SRAM_cell1_dummy_R_64x8m81_1 a_23341_1594# ypass_gate_64x8m81_0_0/bb 018SRAM_cell1_dummy_R_64x8m81_1/a_246_342#
+ 018SRAM_cell1_dummy_R_64x8m81_8/a_126_298# 018SRAM_cell1_dummy_R_64x8m81_1/m3_n36_330#
+ ypass_gate_64x8m81_0_0/b 018SRAM_cell1_dummy_R_64x8m81_8/w_n68_622# vss x018SRAM_cell1_dummy_R_64x8m81
Xnmos_5p04310589983256_64x8m81_0 pmos_5p04310589983254_64x8m81_0/D ypass_gate_64x8m81_0_0/d
+ vss ypass_gate_64x8m81_0_0/d vss nmos_5p04310589983256_64x8m81
X018SRAM_cell1_dummy_R_64x8m81_2 DWL ypass_gate_64x8m81_0_0/bb vss 018SRAM_cell1_64x8m81_1/w_n68_622#
+ DWL ypass_gate_64x8m81_0_0/b 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_R_64x8m81
X018SRAM_cell1_2x_64x8m81_0 018SRAM_cell1_2x_64x8m81_0/018SRAM_cell1_64x8m81_1/m3_n36_330#
+ 018SRAM_cell1_2x_64x8m81_0/018SRAM_cell1_64x8m81_0/m3_n36_330# vss 018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_64x8m81_1/a_444_n42# vss 018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_64x8m81_1/a_36_n42#
+ a_n257_1594# a_n257_1594# 018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ vss x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_dummy_R_64x8m81_3 a_23341_1594# ypass_gate_64x8m81_0_0/bb 018SRAM_cell1_dummy_R_64x8m81_3/a_246_342#
+ 018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_dummy_R_64x8m81_3/m3_n36_330# ypass_gate_64x8m81_0_0/b
+ 018SRAM_cell1_64x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_R_64x8m81
.ends

.subckt rcol4_64_64x8m81 pcb[6] pcb[7] pcb[4] vdd WEN[4] WEN[7] pcb[5] WEN[5] WEN[6]
+ WL[6] WL[5] ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] DWL tblhl GWEN
+ ypass[0] WL[0] WL[2] WL[3] WL[4] WL[7] WL[1] ypass[7] din[4] din[7] q[5] q[6] q[7]
+ din[5] din[6] q[4] a_17474_27175# men col_64a_64x8m81_0/WL[0] rdummy_64x4_64x8m81_0/pcb
+ a_17474_27950# col_64a_64x8m81_0/WL[1] col_64a_64x8m81_0/WL[2] col_64a_64x8m81_0/WL[3]
+ col_64a_64x8m81_0/WL[4] col_64a_64x8m81_0/WL[5] col_64a_64x8m81_0/WL[6] col_64a_64x8m81_0/WL[7]
+ a_6674_27175# rdummy_64x4_64x8m81_0/DWL a_6674_27950# a_17234_27175# a_17234_27950#
+ saout_R_m2_64x8m81_1/WEN rdummy_64x4_64x8m81_0/a_23395_52# a_6434_27175# a_6434_27950#
+ saout_m2_64x8m81_1/mux821_64x8m81_0/a_656_7735# m3_n1_30537# rdummy_64x4_64x8m81_0/a_23341_1594#
+ rdummy_64x4_64x8m81_0/VSS saout_R_m2_64x8m81_1/pcb saout_m2_64x8m81_1/sa_64x8m81_0/pcb
+ saout_R_m2_64x8m81_0/sa_64x8m81_0/pcb saout_m2_64x8m81_0/pcb GWE VSS VDD
Xdcap_103_novia_64x8m81_0[0] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[1] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[2] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[3] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[4] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[5] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[6] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[7] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[8] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[9] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[10] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[11] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[12] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[13] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[14] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[15] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[16] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[17] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[18] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[19] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[20] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[21] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[22] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[23] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[24] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[25] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[26] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[27] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[28] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[29] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[30] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[31] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[32] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[33] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[34] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[35] VDD VDD VSS dcap_103_novia_64x8m81
Xsaout_R_m2_64x8m81_0 saout_R_m2_64x8m81_0/pcb saout_R_m2_64x8m81_0/datain saout_R_m2_64x8m81_0/WEN
+ ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7] men ypass[0] GWEN
+ col_64a_64x8m81_0/BL saout_R_m2_64x8m81_0/q col_64a_64x8m81_0/BL saout_R_m2_64x8m81_0/sa_64x8m81_0/wep
+ saout_R_m2_64x8m81_0/outbuf_oe_64x8m81_0/a_4913_n316# GWE saout_R_m2_64x8m81_0/bb[2]
+ col_64a_64x8m81_0/BL1B col_64a_64x8m81_0/BL ypass[7] saout_R_m2_64x8m81_0/bb[0]
+ saout_R_m2_64x8m81_0/sacntl_2_64x8m81_0/a_4560_1922# saout_m2_64x8m81_1/mux821_64x8m81_0/a_656_7735#
+ col_64a_64x8m81_0/BL1B GWEN a_6900_27175# a_6674_27175# col_64a_64x8m81_0/BL col_64a_64x8m81_0/BL
+ col_64a_64x8m81_0/BL a_6900_27950# a_6674_27950# col_64a_64x8m81_0/BL1B col_64a_64x8m81_0/BL1B
+ saout_R_m2_64x8m81_0/bb[4] men col_64a_64x8m81_0/BL ypass[0] saout_R_m2_64x8m81_0/bb[6]
+ ypass[2] ypass[1] saout_R_m2_64x8m81_0/wen_wm1_64x8m81_0/wen ypass[5] VDD col_64a_64x8m81_0/BL
+ ypass[6] saout_R_m2_64x8m81_0/sa_64x8m81_0/pcb saout_R_m2_64x8m81_0/sacntl_2_64x8m81_0/a_4718_983#
+ saout_R_m2_64x8m81_0/mux821_64x8m81_0/ypass_gate_64x8m81_4/b ypass[3] ypass[4] VSS
+ VDD VDD VDD saout_R_m2_64x8m81
Xcol_64a_64x8m81_0 col_64a_64x8m81_0/WL[0] col_64a_64x8m81_0/WL[6] col_64a_64x8m81_0/WL[4]
+ col_64a_64x8m81_0/WL[3] col_64a_64x8m81_0/WL[7] col_64a_64x8m81_0/WL[1] saout_R_m2_64x8m81_1/bb[2]
+ col_64a_64x8m81_0/b[5] saout_m2_64x8m81_1/bb[5] col_64a_64x8m81_0/b[1] saout_R_m2_64x8m81_0/bb[0]
+ saout_R_m2_64x8m81_0/bb[6] col_64a_64x8m81_0/b[7] saout_R_m2_64x8m81_1/bb[6] saout_m2_64x8m81_0/bb[3]
+ col_64a_64x8m81_0/WL[5] saout_m2_64x8m81_0/bb[5] saout_m2_64x8m81_0/bb[1] col_64a_64x8m81_0/b[3]
+ saout_R_m2_64x8m81_0/bb[2] saout_m2_64x8m81_0/b[4] col_64a_64x8m81_0/b[6] saout_R_m2_64x8m81_0/bb[4]
+ col_64a_64x8m81_0/b[4] saout_R_m2_64x8m81_1/bb[4] saout_R_m2_64x8m81_1/bb[0] col_64a_64x8m81_0/WL[2]
+ saout_m2_64x8m81_1/bb[3] saout_m2_64x8m81_1/bb[7] col_64a_64x8m81_0/BL col_64a_64x8m81_0/bb[7]
+ col_64a_64x8m81_0/BL1B saout_m2_64x8m81_1/bb[1] VSS col_64a_64x8m81_0/b[0] VDD col_64a_64x8m81
Xsaout_R_m2_64x8m81_1 saout_R_m2_64x8m81_1/pcb saout_R_m2_64x8m81_1/datain saout_R_m2_64x8m81_1/WEN
+ ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7] men ypass[0] GWEN
+ col_64a_64x8m81_0/BL saout_R_m2_64x8m81_1/q col_64a_64x8m81_0/BL saout_R_m2_64x8m81_1/sa_64x8m81_0/wep
+ saout_R_m2_64x8m81_1/outbuf_oe_64x8m81_0/a_4913_n316# GWE saout_R_m2_64x8m81_1/bb[2]
+ col_64a_64x8m81_0/BL1B col_64a_64x8m81_0/BL ypass[7] saout_R_m2_64x8m81_1/bb[0]
+ saout_R_m2_64x8m81_1/sacntl_2_64x8m81_0/a_4560_1922# saout_m2_64x8m81_1/mux821_64x8m81_0/a_656_7735#
+ col_64a_64x8m81_0/BL1B GWEN a_17700_27175# a_17474_27175# col_64a_64x8m81_0/BL col_64a_64x8m81_0/BL
+ col_64a_64x8m81_0/BL a_17700_27950# a_17474_27950# col_64a_64x8m81_0/BL1B col_64a_64x8m81_0/BL1B
+ saout_R_m2_64x8m81_1/bb[4] men col_64a_64x8m81_0/BL ypass[0] saout_R_m2_64x8m81_1/bb[6]
+ ypass[2] ypass[1] saout_R_m2_64x8m81_1/wen_wm1_64x8m81_0/wen ypass[5] VDD col_64a_64x8m81_0/BL
+ ypass[6] saout_R_m2_64x8m81_1/pcb saout_R_m2_64x8m81_1/sacntl_2_64x8m81_0/a_4718_983#
+ saout_R_m2_64x8m81_1/mux821_64x8m81_0/ypass_gate_64x8m81_4/b ypass[3] ypass[4] VSS
+ VDD VDD VDD saout_R_m2_64x8m81
Xsaout_m2_64x8m81_0 saout_m2_64x8m81_0/pcb saout_m2_64x8m81_0/datain saout_m2_64x8m81_0/WEN
+ ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7] men ypass[0] GWEN
+ saout_m2_64x8m81_0/bb[5] col_64a_64x8m81_0/b[6] col_64a_64x8m81_0/BL1B saout_m2_64x8m81_0/q
+ a_17009_27175# a_17234_27175# saout_m2_64x8m81_0/sa_64x8m81_0/wep a_17009_27950#
+ a_17234_27950# VSS GWE saout_m2_64x8m81_0/mux821_64x8m81_0/a_4992_424# saout_m2_64x8m81_0/b[4]
+ col_64a_64x8m81_0/BL col_64a_64x8m81_0/bb[7] VSS saout_m2_64x8m81_1/mux821_64x8m81_0/a_656_7735#
+ GWEN ypass[7] col_64a_64x8m81_0/b[7] col_64a_64x8m81_0/b[5] col_64a_64x8m81_0/b[1]
+ col_64a_64x8m81_0/b[4] col_64a_64x8m81_0/BL1B col_64a_64x8m81_0/BL1B saout_m2_64x8m81_0/bb[3]
+ col_64a_64x8m81_0/b[3] saout_m2_64x8m81_0/mux821_64x8m81_0/ypass_gate_a_64x8m81_0/a_n80_n10#
+ ypass[0] saout_m2_64x8m81_0/bb[1] ypass[2] ypass[1] VDD col_64a_64x8m81_0/b[0] saout_m2_64x8m81_0/pcb
+ VSS men ypass[5] VDD ypass[3] ypass[4] col_64a_64x8m81_0/BL1B ypass[6] VSS VDD VDD
+ saout_m2_64x8m81
Xsaout_m2_64x8m81_1 saout_m2_64x8m81_1/pcb saout_m2_64x8m81_1/datain saout_m2_64x8m81_1/WEN
+ ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7] men ypass[0] GWEN
+ saout_m2_64x8m81_1/bb[5] col_64a_64x8m81_0/BL col_64a_64x8m81_0/BL1B saout_m2_64x8m81_1/q
+ a_6209_27175# a_6434_27175# saout_m2_64x8m81_1/sa_64x8m81_0/wep a_6209_27950# a_6434_27950#
+ VSS GWE saout_m2_64x8m81_1/mux821_64x8m81_0/a_4992_424# col_64a_64x8m81_0/BL1B col_64a_64x8m81_0/BL
+ saout_m2_64x8m81_1/bb[7] saout_m2_64x8m81_1/sacntl_2_64x8m81_0/a_4560_1922# saout_m2_64x8m81_1/mux821_64x8m81_0/a_656_7735#
+ GWEN ypass[7] col_64a_64x8m81_0/BL col_64a_64x8m81_0/BL col_64a_64x8m81_0/BL col_64a_64x8m81_0/BL
+ col_64a_64x8m81_0/BL1B col_64a_64x8m81_0/BL1B saout_m2_64x8m81_1/bb[3] col_64a_64x8m81_0/BL
+ saout_m2_64x8m81_1/mux821_64x8m81_0/ypass_gate_a_64x8m81_0/a_n80_n10# ypass[0] saout_m2_64x8m81_1/bb[1]
+ ypass[2] ypass[1] VDD col_64a_64x8m81_0/BL saout_m2_64x8m81_1/sa_64x8m81_0/pcb saout_m2_64x8m81_1/sacntl_2_64x8m81_0/a_4718_983#
+ men ypass[5] VDD ypass[3] ypass[4] saout_m2_64x8m81_1/mux821_64x8m81_0/ypass_gate_a_64x8m81_0/b
+ ypass[6] VSS VDD VDD saout_m2_64x8m81
Xrdummy_64x4_64x8m81_0 tblhl rdummy_64x4_64x8m81_0/pcb col_64a_64x8m81_0/BL1B ypass[1]
+ saout_m2_64x8m81_0/bb[1] col_64a_64x8m81_0/BL1B VSS col_64a_64x8m81_0/BL1B col_64a_64x8m81_0/WL[4]
+ saout_R_m2_64x8m81_1/bb[2] col_64a_64x8m81_0/BL rdummy_64x4_64x8m81_0/ypass_gate_64x8m81_0_0/d
+ col_64a_64x8m81_0/WL[2] col_64a_64x8m81_0/BL col_64a_64x8m81_0/BL1B col_64a_64x8m81_0/BL
+ saout_R_m2_64x8m81_1/bb[0] col_64a_64x8m81_0/BL VDD col_64a_64x8m81_0/BL1B col_64a_64x8m81_0/WL[0]
+ ypass[6] col_64a_64x8m81_0/b[0] col_64a_64x8m81_0/b[0] VSS VSS col_64a_64x8m81_0/b[1]
+ col_64a_64x8m81_0/BL1B col_64a_64x8m81_0/WL[6] col_64a_64x8m81_0/b[1] col_64a_64x8m81_0/WL[1]
+ col_64a_64x8m81_0/BL1B col_64a_64x8m81_0/BL col_64a_64x8m81_0/WL[5] col_64a_64x8m81_0/BL
+ col_64a_64x8m81_0/BL col_64a_64x8m81_0/b[3] col_64a_64x8m81_0/BL col_64a_64x8m81_0/WL[7]
+ col_64a_64x8m81_0/BL col_64a_64x8m81_0/WL[2] saout_m2_64x8m81_0/bb[3] col_64a_64x8m81_0/b[5]
+ col_64a_64x8m81_0/WL[3] VSS col_64a_64x8m81_0/b[4] saout_m2_64x8m81_1/bb[7] col_64a_64x8m81_0/WL[1]
+ saout_m2_64x8m81_1/bb[1] col_64a_64x8m81_0/b[6] col_64a_64x8m81_0/BL col_64a_64x8m81_0/BL
+ col_64a_64x8m81_0/b[7] col_64a_64x8m81_0/BL saout_m2_64x8m81_0/bb[5] saout_m2_64x8m81_0/bb[3]
+ VSS col_64a_64x8m81_0/BL rdummy_64x4_64x8m81_0/DWL col_64a_64x8m81_0/BL col_64a_64x8m81_0/BL1B
+ col_64a_64x8m81_0/BL1B col_64a_64x8m81_0/b[3] col_64a_64x8m81_0/BL1B col_64a_64x8m81_0/BL1B
+ col_64a_64x8m81_0/BL rdummy_64x4_64x8m81_0/a_23395_52# col_64a_64x8m81_0/BL col_64a_64x8m81_0/b[5]
+ saout_R_m2_64x8m81_1/bb[6] saout_m2_64x8m81_0/b[4] saout_m2_64x8m81_0/bb[5] col_64a_64x8m81_0/b[4]
+ VSS col_64a_64x8m81_0/BL saout_R_m2_64x8m81_1/bb[4] ypass[0] col_64a_64x8m81_0/b[6]
+ saout_m2_64x8m81_1/bb[3] col_64a_64x8m81_0/BL1B col_64a_64x8m81_0/b[7] saout_m2_64x8m81_1/bb[1]
+ col_64a_64x8m81_0/BL1B col_64a_64x8m81_0/BL col_64a_64x8m81_0/BL1B col_64a_64x8m81_0/BL
+ VDD saout_R_m2_64x8m81_1/bb[2] col_64a_64x8m81_0/BL1B ypass[5] saout_m2_64x8m81_0/b[4]
+ VSS col_64a_64x8m81_0/BL col_64a_64x8m81_0/WL[3] col_64a_64x8m81_0/BL1B saout_R_m2_64x8m81_1/bb[0]
+ col_64a_64x8m81_0/WL[6] saout_R_m2_64x8m81_0/bb[2] saout_m2_64x8m81_1/bb[5] saout_R_m2_64x8m81_0/bb[6]
+ col_64a_64x8m81_0/WL[4] col_64a_64x8m81_0/BL1B col_64a_64x8m81_0/BL1B saout_R_m2_64x8m81_0/bb[4]
+ col_64a_64x8m81_0/BL col_64a_64x8m81_0/BL saout_R_m2_64x8m81_0/bb[0] col_64a_64x8m81_0/bb[7]
+ col_64a_64x8m81_0/BL1B col_64a_64x8m81_0/BL1B col_64a_64x8m81_0/BL VDD rdummy_64x4_64x8m81_0/a_23341_1594#
+ col_64a_64x8m81_0/BL col_64a_64x8m81_0/BL1B col_64a_64x8m81_0/BL col_64a_64x8m81_0/BL1B
+ saout_R_m2_64x8m81_0/bb[2] col_64a_64x8m81_0/BL col_64a_64x8m81_0/BL1B col_64a_64x8m81_0/BL
+ col_64a_64x8m81_0/BL col_64a_64x8m81_0/BL VDD saout_R_m2_64x8m81_0/bb[0] col_64a_64x8m81_0/bb[7]
+ ypass[2] col_64a_64x8m81_0/BL col_64a_64x8m81_0/BL col_64a_64x8m81_0/BL VDD col_64a_64x8m81_0/BL
+ rdummy_64x4_64x8m81_0/ypass_gate_64x8m81_0_0/d col_64a_64x8m81_0/BL1B col_64a_64x8m81_0/BL
+ ypass[4] col_64a_64x8m81_0/BL col_64a_64x8m81_0/BL col_64a_64x8m81_0/BL col_64a_64x8m81_0/BL
+ col_64a_64x8m81_0/BL VDD col_64a_64x8m81_0/BL1B col_64a_64x8m81_0/BL col_64a_64x8m81_0/BL
+ col_64a_64x8m81_0/BL VSS col_64a_64x8m81_0/BL col_64a_64x8m81_0/BL col_64a_64x8m81_0/WL[7]
+ rdummy_64x4_64x8m81_0/VSS col_64a_64x8m81_0/BL saout_m2_64x8m81_0/bb[1] VDD col_64a_64x8m81_0/BL1B
+ col_64a_64x8m81_0/WL[5] ypass[3] VSS col_64a_64x8m81_0/WL[0] saout_m2_64x8m81_1/bb[3]
+ saout_R_m2_64x8m81_0/bb[6] VDD m3_n1_30537# col_64a_64x8m81_0/BL saout_R_m2_64x8m81_0/bb[4]
+ col_64a_64x8m81_0/BL col_64a_64x8m81_0/BL1B saout_m2_64x8m81_1/bb[7] col_64a_64x8m81_0/BL1B
+ VDD col_64a_64x8m81_0/BL1B col_64a_64x8m81_0/BL1B saout_m2_64x8m81_1/bb[5] VDD saout_R_m2_64x8m81_1/bb[6]
+ VSS col_64a_64x8m81_0/BL ypass[7] col_64a_64x8m81_0/BL saout_R_m2_64x8m81_1/bb[4]
+ VSS col_64a_64x8m81_0/BL rdummy_64x4_64x8m81
.ends

.subckt pmos_5p043105899832101_64x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=6.59u l=0.6u
.ends

.subckt pmoscap_W2_5_477_R270_64x8m81 m3_489_n1# m3_1409_n1# w_n60_n407# a_81_507#
X0 a_81_507# a_49_1969# a_81_507# w_n60_n407# pmos_3p3 w=5.495u l=3.94u
X1 a_81_507# a_49_1969# a_81_507# w_n60_n407# pmos_3p3 w=5.495u l=3.94u
.ends

.subckt pmos_5p043105899832111_64x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.59u l=0.6u
.ends

.subckt pmos_5p043105899832106_64x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=3.3u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=3.3u l=0.6u
.ends

.subckt pmos_1p2$$49271852_R270_64x8m81 w_n296_n137# pmos_5p043105899832106_64x8m81_0/S
+ pmos_5p043105899832106_64x8m81_0/D a_193_n71# a_n31_n71#
Xpmos_5p043105899832106_64x8m81_0 w_n296_n137# pmos_5p043105899832106_64x8m81_0/D
+ a_n31_n71# pmos_5p043105899832106_64x8m81_0/S a_193_n71# pmos_5p043105899832106_64x8m81
.ends

.subckt nmos_5p043105899832109_64x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=5u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=5u l=0.6u
.ends

.subckt nmos_5p043105899832110_64x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=3.3u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=3.3u l=0.6u
.ends

.subckt pmos_5p043105899832104_64x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.62u l=0.6u
.ends

.subckt pmos_5p043105899832108_64x8m81 w_n208_n120# D a_0_n44# S a_448_n44# a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=10u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=10u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=10u l=0.6u
.ends

.subckt pmos_1p2$$49270828_R270_64x8m81 w_n296_n137# pmos_5p043105899832108_64x8m81_0/S
+ a_193_n71# pmos_5p043105899832108_64x8m81_0/D a_n31_n71# a_417_n71#
Xpmos_5p043105899832108_64x8m81_0 w_n296_n137# pmos_5p043105899832108_64x8m81_0/D
+ a_n31_n71# pmos_5p043105899832108_64x8m81_0/S a_417_n71# a_193_n71# pmos_5p043105899832108_64x8m81
.ends

.subckt nmos_5p043105899832107_64x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=0.66u l=0.6u
.ends

.subckt pmos_5p043105899832105_64x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=5.5u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=5.5u l=0.6u
.ends

.subckt pmos_1p2$$49272876_R270_64x8m81 w_n296_n137# pmos_5p043105899832105_64x8m81_0/S
+ pmos_5p043105899832105_64x8m81_0/D a_n31_n71# a_193_n71#
Xpmos_5p043105899832105_64x8m81_0 w_n296_n137# pmos_5p043105899832105_64x8m81_0/D
+ a_n31_n71# pmos_5p043105899832105_64x8m81_0/S a_193_n71# pmos_5p043105899832105_64x8m81
.ends

.subckt nmos_1p2$$49277996_R270_64x8m81 nmos_5p04310589983249_64x8m81_0/S a_n31_n71#
+ nmos_5p04310589983249_64x8m81_0/D VSUBS
Xnmos_5p04310589983249_64x8m81_0 nmos_5p04310589983249_64x8m81_0/D a_n31_n71# nmos_5p04310589983249_64x8m81_0/S
+ VSUBS nmos_5p04310589983249_64x8m81
.ends

.subckt xdec_64x8m81 xc xb xa RWL LWL m2_16621_n223# m2_17754_n223# m2_11825_n223#
+ m2_12202_n223# m2_12958_n223# m2_15487_n223# m2_12580_n223# m2_15110_n223# m2_11069_n223#
+ m2_15865_n223# m2_16243_n223# men m2_10314_n223# vss m2_16998_n223# m2_17376_n223#
+ m2_11447_n223# m2_10691_n223# vdd
Xpmos_5p043105899832111_64x8m81_0 vdd vdd pmos_5p043105899832104_64x8m81_2/S pmos_5p043105899832111_64x8m81_0/S
+ pmos_5p043105899832111_64x8m81
Xpmos_1p2$$49271852_R270_64x8m81_0 vdd nmos_5p043105899832110_64x8m81_0/S men pmos_5p043105899832104_64x8m81_2/S
+ pmos_5p043105899832104_64x8m81_2/S pmos_1p2$$49271852_R270_64x8m81
Xnmos_5p043105899832109_64x8m81_0 LWL pmos_1p2$$49272876_R270_64x8m81_1/pmos_5p043105899832105_64x8m81_0/D
+ vss pmos_1p2$$49272876_R270_64x8m81_1/pmos_5p043105899832105_64x8m81_0/D vss nmos_5p043105899832109_64x8m81
Xnmos_5p043105899832109_64x8m81_1 RWL pmos_1p2$$49272876_R270_64x8m81_0/pmos_5p043105899832105_64x8m81_0/D
+ vss pmos_1p2$$49272876_R270_64x8m81_0/pmos_5p043105899832105_64x8m81_0/D vss nmos_5p043105899832109_64x8m81
Xnmos_5p043105899832110_64x8m81_0 men pmos_5p043105899832111_64x8m81_0/S nmos_5p043105899832110_64x8m81_0/S
+ pmos_5p043105899832111_64x8m81_0/S vss nmos_5p043105899832110_64x8m81
Xpmos_5p043105899832104_64x8m81_0 vdd pmos_5p043105899832104_64x8m81_2/S xb vdd pmos_5p043105899832104_64x8m81
Xpmos_5p043105899832108_64x8m81_0 vdd vdd pmos_1p2$$49272876_R270_64x8m81_0/pmos_5p043105899832105_64x8m81_0/D
+ RWL pmos_1p2$$49272876_R270_64x8m81_0/pmos_5p043105899832105_64x8m81_0/D pmos_1p2$$49272876_R270_64x8m81_0/pmos_5p043105899832105_64x8m81_0/D
+ pmos_5p043105899832108_64x8m81
Xpmos_5p043105899832104_64x8m81_1 vdd vdd xc pmos_5p043105899832104_64x8m81_2/S pmos_5p043105899832104_64x8m81
Xpmos_5p043105899832104_64x8m81_2 vdd vdd xa pmos_5p043105899832104_64x8m81_2/S pmos_5p043105899832104_64x8m81
Xpmos_1p2$$49270828_R270_64x8m81_0 vdd LWL pmos_1p2$$49272876_R270_64x8m81_1/pmos_5p043105899832105_64x8m81_0/D
+ vdd pmos_1p2$$49272876_R270_64x8m81_1/pmos_5p043105899832105_64x8m81_0/D pmos_1p2$$49272876_R270_64x8m81_1/pmos_5p043105899832105_64x8m81_0/D
+ pmos_1p2$$49270828_R270_64x8m81
Xnmos_5p043105899832107_64x8m81_0 vss pmos_5p043105899832104_64x8m81_2/S pmos_5p043105899832111_64x8m81_0/S
+ vss nmos_5p043105899832107_64x8m81
Xpmos_1p2$$49272876_R270_64x8m81_0 vdd vdd pmos_1p2$$49272876_R270_64x8m81_0/pmos_5p043105899832105_64x8m81_0/D
+ nmos_5p043105899832110_64x8m81_0/S nmos_5p043105899832110_64x8m81_0/S pmos_1p2$$49272876_R270_64x8m81
Xpmos_1p2$$49272876_R270_64x8m81_1 vdd vdd pmos_1p2$$49272876_R270_64x8m81_1/pmos_5p043105899832105_64x8m81_0/D
+ nmos_5p043105899832110_64x8m81_0/S nmos_5p043105899832110_64x8m81_0/S pmos_1p2$$49272876_R270_64x8m81
Xnmos_1p2$$49277996_R270_64x8m81_0 nmos_5p043105899832110_64x8m81_0/S pmos_5p043105899832104_64x8m81_2/S
+ vss vss nmos_1p2$$49277996_R270_64x8m81
X0 a_13291_624# xb a_13291_400# vss nmos_3p3 w=3.15u l=0.6u
X1 vss xc a_13291_624# vss nmos_3p3 w=3.15u l=0.6u
X2 a_13291_400# xa pmos_5p043105899832104_64x8m81_2/S vss nmos_3p3 w=3.15u l=0.6u
X3 vss nmos_5p043105899832110_64x8m81_0/S pmos_1p2$$49272876_R270_64x8m81_0/pmos_5p043105899832105_64x8m81_0/D vss nmos_3p3 w=5u l=0.6u
X4 vss nmos_5p043105899832110_64x8m81_0/S pmos_1p2$$49272876_R270_64x8m81_1/pmos_5p043105899832105_64x8m81_0/D vss nmos_3p3 w=5u l=0.6u
.ends

.subckt xdec8_64x8m81 xb xa[4] xa[6] xa[7] xa[1] RWL[0] LWL[5] LWL[4] LWL[2] RWL[4]
+ RWL[1] RWL[7] RWL[6] LWL[1] LWL[7] RWL[3] xdec_64x8m81_3/RWL xa[3] xa[0] xdec_64x8m81_7/m2_17754_n223#
+ xdec_64x8m81_7/m2_11825_n223# xdec_64x8m81_7/m2_12202_n223# xdec_64x8m81_7/m2_10314_n223#
+ RWL[5] xdec_64x8m81_7/m2_11069_n223# xdec_64x8m81_7/m2_17376_n223# xdec_64x8m81_7/m2_12958_n223#
+ xdec_64x8m81_7/m2_15110_n223# LWL[3] xc xdec_64x8m81_7/m2_15487_n223# xa[5] RWL[2]
+ xa[2] xdec_64x8m81_7/m2_15865_n223# LWL[0] xdec_64x8m81_7/m2_11447_n223# xdec_64x8m81_7/m2_16243_n223#
+ xdec_64x8m81_7/m2_12580_n223# LWL[6] xdec_64x8m81_7/m2_16621_n223# xdec_64x8m81_7/m2_10691_n223#
+ vdd xdec_64x8m81_7/m2_16998_n223# vss men
Xxdec_64x8m81_0 xc xb xa[6] RWL[6] LWL[6] xdec_64x8m81_7/m2_16621_n223# xdec_64x8m81_7/m2_17754_n223#
+ xdec_64x8m81_7/m2_11825_n223# xdec_64x8m81_7/m2_12202_n223# xdec_64x8m81_7/m2_12958_n223#
+ xdec_64x8m81_7/m2_15487_n223# xdec_64x8m81_7/m2_12580_n223# xdec_64x8m81_7/m2_15110_n223#
+ xdec_64x8m81_7/m2_11069_n223# xdec_64x8m81_7/m2_15865_n223# xdec_64x8m81_7/m2_16243_n223#
+ men xdec_64x8m81_7/m2_10314_n223# vss xdec_64x8m81_7/m2_16998_n223# xdec_64x8m81_7/m2_17376_n223#
+ xdec_64x8m81_7/m2_11447_n223# xdec_64x8m81_7/m2_10691_n223# vdd xdec_64x8m81
Xxdec_64x8m81_1 xc xb xa[4] RWL[4] LWL[4] xdec_64x8m81_7/m2_16621_n223# xdec_64x8m81_7/m2_17754_n223#
+ xdec_64x8m81_7/m2_11825_n223# xdec_64x8m81_7/m2_12202_n223# xdec_64x8m81_7/m2_12958_n223#
+ xdec_64x8m81_7/m2_15487_n223# xdec_64x8m81_7/m2_12580_n223# xdec_64x8m81_7/m2_15110_n223#
+ xdec_64x8m81_7/m2_11069_n223# xdec_64x8m81_7/m2_15865_n223# xdec_64x8m81_7/m2_16243_n223#
+ men xdec_64x8m81_7/m2_10314_n223# vss xdec_64x8m81_7/m2_16998_n223# xdec_64x8m81_7/m2_17376_n223#
+ xdec_64x8m81_7/m2_11447_n223# xdec_64x8m81_7/m2_10691_n223# vdd xdec_64x8m81
Xxdec_64x8m81_2 xc xb xa[2] RWL[2] LWL[2] xdec_64x8m81_7/m2_16621_n223# xdec_64x8m81_7/m2_17754_n223#
+ xdec_64x8m81_7/m2_11825_n223# xdec_64x8m81_7/m2_12202_n223# xdec_64x8m81_7/m2_12958_n223#
+ xdec_64x8m81_7/m2_15487_n223# xdec_64x8m81_7/m2_12580_n223# xdec_64x8m81_7/m2_15110_n223#
+ xdec_64x8m81_7/m2_11069_n223# xdec_64x8m81_7/m2_15865_n223# xdec_64x8m81_7/m2_16243_n223#
+ men xdec_64x8m81_7/m2_10314_n223# vss xdec_64x8m81_7/m2_16998_n223# xdec_64x8m81_7/m2_17376_n223#
+ xdec_64x8m81_7/m2_11447_n223# xdec_64x8m81_7/m2_10691_n223# vdd xdec_64x8m81
Xxdec_64x8m81_3 xc xb xa[0] xdec_64x8m81_3/RWL LWL[0] xdec_64x8m81_7/m2_16621_n223#
+ xdec_64x8m81_7/m2_17754_n223# xdec_64x8m81_7/m2_11825_n223# xdec_64x8m81_7/m2_12202_n223#
+ xdec_64x8m81_7/m2_12958_n223# xdec_64x8m81_7/m2_15487_n223# xdec_64x8m81_7/m2_12580_n223#
+ xdec_64x8m81_7/m2_15110_n223# xdec_64x8m81_7/m2_11069_n223# xdec_64x8m81_7/m2_15865_n223#
+ xdec_64x8m81_7/m2_16243_n223# men xdec_64x8m81_7/m2_10314_n223# vss xdec_64x8m81_7/m2_16998_n223#
+ xdec_64x8m81_7/m2_17376_n223# xdec_64x8m81_7/m2_11447_n223# xdec_64x8m81_7/m2_10691_n223#
+ vdd xdec_64x8m81
Xxdec_64x8m81_4 xc xb xa[7] RWL[7] LWL[7] xdec_64x8m81_7/m2_16621_n223# xdec_64x8m81_7/m2_17754_n223#
+ xdec_64x8m81_7/m2_11825_n223# xdec_64x8m81_7/m2_12202_n223# xdec_64x8m81_7/m2_12958_n223#
+ xdec_64x8m81_7/m2_15487_n223# xdec_64x8m81_7/m2_12580_n223# xdec_64x8m81_7/m2_15110_n223#
+ xdec_64x8m81_7/m2_11069_n223# xdec_64x8m81_7/m2_15865_n223# xdec_64x8m81_7/m2_16243_n223#
+ men xdec_64x8m81_7/m2_10314_n223# vss xdec_64x8m81_7/m2_16998_n223# xdec_64x8m81_7/m2_17376_n223#
+ xdec_64x8m81_7/m2_11447_n223# xdec_64x8m81_7/m2_10691_n223# vdd xdec_64x8m81
Xxdec_64x8m81_5 xc xb xa[5] RWL[5] LWL[5] xdec_64x8m81_7/m2_16621_n223# xdec_64x8m81_7/m2_17754_n223#
+ xdec_64x8m81_7/m2_11825_n223# xdec_64x8m81_7/m2_12202_n223# xdec_64x8m81_7/m2_12958_n223#
+ xdec_64x8m81_7/m2_15487_n223# xdec_64x8m81_7/m2_12580_n223# xdec_64x8m81_7/m2_15110_n223#
+ xdec_64x8m81_7/m2_11069_n223# xdec_64x8m81_7/m2_15865_n223# xdec_64x8m81_7/m2_16243_n223#
+ men xdec_64x8m81_7/m2_10314_n223# vss xdec_64x8m81_7/m2_16998_n223# xdec_64x8m81_7/m2_17376_n223#
+ xdec_64x8m81_7/m2_11447_n223# xdec_64x8m81_7/m2_10691_n223# vdd xdec_64x8m81
Xxdec_64x8m81_6 xc xb xa[3] RWL[3] LWL[3] xdec_64x8m81_7/m2_16621_n223# xdec_64x8m81_7/m2_17754_n223#
+ xdec_64x8m81_7/m2_11825_n223# xdec_64x8m81_7/m2_12202_n223# xdec_64x8m81_7/m2_12958_n223#
+ xdec_64x8m81_7/m2_15487_n223# xdec_64x8m81_7/m2_12580_n223# xdec_64x8m81_7/m2_15110_n223#
+ xdec_64x8m81_7/m2_11069_n223# xdec_64x8m81_7/m2_15865_n223# xdec_64x8m81_7/m2_16243_n223#
+ men xdec_64x8m81_7/m2_10314_n223# vss xdec_64x8m81_7/m2_16998_n223# xdec_64x8m81_7/m2_17376_n223#
+ xdec_64x8m81_7/m2_11447_n223# xdec_64x8m81_7/m2_10691_n223# vdd xdec_64x8m81
Xxdec_64x8m81_7 xc xb xa[1] RWL[1] LWL[1] xdec_64x8m81_7/m2_16621_n223# xdec_64x8m81_7/m2_17754_n223#
+ xdec_64x8m81_7/m2_11825_n223# xdec_64x8m81_7/m2_12202_n223# xdec_64x8m81_7/m2_12958_n223#
+ xdec_64x8m81_7/m2_15487_n223# xdec_64x8m81_7/m2_12580_n223# xdec_64x8m81_7/m2_15110_n223#
+ xdec_64x8m81_7/m2_11069_n223# xdec_64x8m81_7/m2_15865_n223# xdec_64x8m81_7/m2_16243_n223#
+ men xdec_64x8m81_7/m2_10314_n223# vss xdec_64x8m81_7/m2_16998_n223# xdec_64x8m81_7/m2_17376_n223#
+ xdec_64x8m81_7/m2_11447_n223# xdec_64x8m81_7/m2_10691_n223# vdd xdec_64x8m81
.ends

.subckt pmos_5p043105899832102_64x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=12.63u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=12.63u l=0.6u
.ends

.subckt pmos_1p2$$204216364_R90_64x8m81 pmos_5p043105899832102_64x8m81_0/S pmos_5p043105899832102_64x8m81_0/D
+ a_193_n71# w_n296_n137# a_n31_n71#
Xpmos_5p043105899832102_64x8m81_0 w_n296_n137# pmos_5p043105899832102_64x8m81_0/D
+ a_n31_n71# pmos_5p043105899832102_64x8m81_0/S a_193_n71# pmos_5p043105899832102_64x8m81
.ends

.subckt nmos_5p04310589983299_64x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=10.11u l=0.6u
.ends

.subckt nmos_1p2$$204213292_R90_64x8m81 nmos_5p04310589983299_64x8m81_0/S a_n31_n71#
+ nmos_5p04310589983299_64x8m81_0/D VSUBS
Xnmos_5p04310589983299_64x8m81_0 nmos_5p04310589983299_64x8m81_0/D a_n31_n71# nmos_5p04310589983299_64x8m81_0/S
+ VSUBS nmos_5p04310589983299_64x8m81
.ends

.subckt nmos_5p043105899832103_64x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=2.64u l=0.6u
.ends

.subckt nmos_5p043105899832100_64x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=6.59u l=0.6u
.ends

.subckt nmos_1p2$$204215_R270_64x8m81 nmos_5p043105899832100_64x8m81_0/S a_n31_n71#
+ nmos_5p043105899832100_64x8m81_0/D VSUBS
Xnmos_5p043105899832100_64x8m81_0 nmos_5p043105899832100_64x8m81_0/D a_n31_n71# nmos_5p043105899832100_64x8m81_0/S
+ VSUBS nmos_5p043105899832100_64x8m81
.ends

.subckt pmoscap_W2_5_R270_64x8m81 w_n60_n407# a_81_507# m3_509_n1#
X0 a_81_507# M1_POLY2$$2043_R270_64x8m81_0/VSUBS a_81_507# w_n60_n407# pmos_3p3 w=5.495u l=3.94u
.ends

.subckt pmos_1p2$$204217388_R90_64x8m81 pmos_5p043105899832101_64x8m81_0/S w_n295_n137#
+ pmos_5p043105899832101_64x8m81_0/D a_n31_n71#
Xpmos_5p043105899832101_64x8m81_0 w_n295_n137# pmos_5p043105899832101_64x8m81_0/D
+ a_n31_n71# pmos_5p043105899832101_64x8m81_0/S pmos_5p043105899832101_64x8m81
.ends

.subckt xdec8_64_64x8m81 DRWL RWL[6] RWL[1] LWL[6] LWL[7] LWL[2] LWL[3] LWL[4] LWL[5]
+ LWL[0] DLWL xa[7] xa[6] xa[5] xa[4] xa[0] xa[3] xa[2] xa[1] RWL[4] RWL[2] RWL[0]
+ men LWL[1] RWL[7] RWL[5] RWL[3] vss vdd
Xpmos_5p043105899832101_64x8m81_0 vdd pmos_5p043105899832101_64x8m81_0/D vss men pmos_5p043105899832101_64x8m81
Xpmoscap_W2_5_477_R270_64x8m81_0 LWL[7] LWL[6] vdd vdd pmoscap_W2_5_477_R270_64x8m81
Xpmos_5p043105899832101_64x8m81_1 vdd vdd pmos_5p043105899832101_64x8m81_0/D pmos_5p043105899832101_64x8m81_1/S
+ pmos_5p043105899832101_64x8m81
Xpmoscap_W2_5_477_R270_64x8m81_1 LWL[5] LWL[4] vdd vdd pmoscap_W2_5_477_R270_64x8m81
Xxdec8_64x8m81_0 vdd xa[4] xa[6] xa[7] xa[1] RWL[0] LWL[5] LWL[4] LWL[2] RWL[4] RWL[1]
+ RWL[7] RWL[6] LWL[1] LWL[7] RWL[3] RWL[0] xa[3] xa[0] xa[0] vdd vdd vdd RWL[5] vdd
+ xa[1] vdd xa[7] LWL[3] vdd xa[6] xa[5] RWL[2] xa[2] xa[5] LWL[0] vdd xa[4] vdd LWL[6]
+ xa[3] vdd vdd xa[2] vss men xdec8_64x8m81
Xpmoscap_W2_5_477_R270_64x8m81_2 LWL[3] LWL[2] vdd vdd pmoscap_W2_5_477_R270_64x8m81
Xpmoscap_W2_5_477_R270_64x8m81_3 LWL[1] LWL[0] vdd vdd pmoscap_W2_5_477_R270_64x8m81
Xpmoscap_W2_5_477_R270_64x8m81_4 RWL[7] RWL[6] vdd vdd pmoscap_W2_5_477_R270_64x8m81
Xpmoscap_W2_5_477_R270_64x8m81_5 RWL[5] RWL[4] vdd vdd pmoscap_W2_5_477_R270_64x8m81
Xpmoscap_W2_5_477_R270_64x8m81_6 RWL[3] RWL[2] vdd vdd pmoscap_W2_5_477_R270_64x8m81
Xpmoscap_W2_5_477_R270_64x8m81_7 RWL[1] RWL[0] vdd vdd pmoscap_W2_5_477_R270_64x8m81
Xpmos_1p2$$204216364_R90_64x8m81_0 vdd DRWL pmos_5p043105899832101_64x8m81_1/S vdd
+ pmos_5p043105899832101_64x8m81_1/S pmos_1p2$$204216364_R90_64x8m81
Xnmos_1p2$$204213292_R90_64x8m81_0 DLWL nmos_5p043105899832103_64x8m81_1/S vss vss
+ nmos_1p2$$204213292_R90_64x8m81
Xpmos_1p2$$204216364_R90_64x8m81_1 vdd DLWL nmos_5p043105899832103_64x8m81_1/S vdd
+ nmos_5p043105899832103_64x8m81_1/S pmos_1p2$$204216364_R90_64x8m81
Xnmos_5p043105899832103_64x8m81_0 vss pmos_5p043105899832101_64x8m81_0/D pmos_5p043105899832101_64x8m81_1/S
+ vss nmos_5p043105899832103_64x8m81
Xnmos_5p043105899832103_64x8m81_1 vss pmos_5p043105899832101_64x8m81_0/D nmos_5p043105899832103_64x8m81_1/S
+ vss nmos_5p043105899832103_64x8m81
Xnmos_1p2$$204215_R270_64x8m81_0 pmos_5p043105899832101_64x8m81_0/D vdd men vss nmos_1p2$$204215_R270_64x8m81
Xpmoscap_W2_5_R270_64x8m81_0 vdd vdd DLWL pmoscap_W2_5_R270_64x8m81
Xpmoscap_W2_5_R270_64x8m81_1 vdd vdd DRWL pmoscap_W2_5_R270_64x8m81
Xpmos_1p2$$204217388_R90_64x8m81_0 nmos_5p043105899832103_64x8m81_1/S vdd vdd pmos_5p043105899832101_64x8m81_0/D
+ pmos_1p2$$204217388_R90_64x8m81
Xnmos_5p04310589983299_64x8m81_0 vss pmos_5p043105899832101_64x8m81_1/S DRWL vss nmos_5p04310589983299_64x8m81
.ends

.subckt x018SRAM_cell1_cutPC_64x8m81 a_n36_52# a_444_n42# a_246_342# a_246_712# m3_n36_330#
+ a_36_n42# w_n68_622# VSUBS
X0 a_126_298# a_n36_52# a_444_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X1 a_36_206# a_n36_52# a_36_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X2 a_246_712# a_126_298# a_36_206# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X3 a_126_298# a_36_206# a_246_712# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X4 a_246_342# a_126_298# a_36_206# VSUBS nmos_6p0 w=0.95u l=0.6u
X5 a_126_298# a_36_206# a_246_342# VSUBS nmos_6p0 w=0.95u l=0.6u
.ends

.subckt new_dummyrow_unit_01_64x8m81 018SRAM_cell1_dummy_64x8m81_12/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_4/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_13/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_5/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_14/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_6/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_15/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_7/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_8/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_0/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_9/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_2/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_1/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_3/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_5/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_4/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_6/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_7/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_0/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_8/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_9/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_10/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_11/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_13/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_12/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_14/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_1/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_15/m2_390_n50#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_10/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_2/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_11/m2_90_n50# VSUBS 018SRAM_cell1_dummy_64x8m81_3/m2_90_n50#
+ 018SRAM_strap1_64x8m81_1/w_n68_622#
X018SRAM_cell1_dummy_64x8m81_10 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_10/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_10/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_11 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_11/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_11/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_12 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_12/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_12/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_13 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_13/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_13/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_14 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_14/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_14/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_15 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_15/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_15/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_0 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_0/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_0/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_1 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_1/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_1/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_2 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_2/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_2/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_3 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_3/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_3/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_5 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_5/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_5/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_4 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_4/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_4/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_6 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_6/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_6/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_7 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_7/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_7/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_8 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_8/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_8/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_9 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_cell1_dummy_64x8m81_9/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_9/m2_390_n50# 018SRAM_strap1_64x8m81_1/w_n68_622#
+ 018SRAM_strap1_64x8m81_1/a_n36_52# 018SRAM_strap1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
.ends

.subckt ldummy_64x4_64x8m81 new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_2/m2_390_n50#
+ 018SRAM_cell1_cutPC_64x8m81_1/m3_n36_330# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_3/m2_390_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_8/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_12/m2_90_n50#
+ 018SRAM_cell1_cutPC_64x8m81_2/m3_n36_330# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_4/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_22/m2_90_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_0/m2_390_n50#
+ 018SRAM_cell1_cutPC_64x8m81_4/a_246_342# 018SRAM_cell1_dummy_64x8m81_4/m2_90_n50#
+ 018SRAM_cell1_cutPC_64x8m81_3/m3_n36_330# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_5/m2_390_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_1/m2_390_n50# 018SRAM_cell1_cutPC_64x8m81_4/m3_n36_330#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_0/m2_90_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_6/m2_390_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_2/m2_390_n50# 018SRAM_cell1_cutPC_64x8m81_5/m3_n36_330#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_7/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_13/m2_90_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_3/m2_390_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_9/m2_90_n50#
+ 018SRAM_cell1_cutPC_64x8m81_6/m3_n36_330# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_8/m2_390_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_4/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_23/m2_90_n50#
+ 018SRAM_cell1_cutPC_64x8m81_5/a_246_342# 018SRAM_cell1_cutPC_64x8m81_7/m3_n36_330#
+ 018SRAM_cell1_cutPC_64x8m81_7/w_n68_622# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_9/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_5/m2_90_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_5/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_1/m2_90_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_6/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_14/m2_90_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_7/m2_390_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_8/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_24/m2_90_n50#
+ 018SRAM_cell1_cutPC_64x8m81_6/a_246_342# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_10/m2_390_n50#
+ 018SRAM_cell1_cutPC_64x8m81_5/w_n68_622# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_9/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_6/m2_90_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_11/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_2/m2_90_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_12/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_10/m2_90_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_0/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_30/m2_390_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_13/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_15/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_25/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_31/m2_390_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_14/m2_390_n50#
+ 018SRAM_cell1_cutPC_64x8m81_7/a_246_342# 018SRAM_cell1_cutPC_64x8m81_4/w_n68_622#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_10/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_7/m2_90_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_15/m2_390_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_11/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_3/m2_90_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_11/m2_90_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_12/m2_390_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_1/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_16/m2_90_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_10/m2_90_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_13/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_26/m2_90_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_14/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_8/m2_90_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_15/m2_390_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_4/m2_90_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_11/m2_90_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_12/m2_90_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_2/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_17/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_27/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_0/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_20/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_9/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_21/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_1/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_5/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_22/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_2/m2_390_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_13/m2_90_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_12/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_23/m2_390_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_3/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_3/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_18/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_24/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_28/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_4/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_5/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_25/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_6/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_6/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_26/m2_390_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_14/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_7/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_19/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_27/m2_390_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_4/m2_90_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_13/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_28/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_29/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_8/m2_390_n50#
+ 018SRAM_cell1_cutPC_64x8m81_0/a_246_342# 018SRAM_cell1_cutPC_64x8m81_7/a_246_712#
+ 018SRAM_cell1_dummy_64x8m81_0/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_10/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_9/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_29/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_7/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_11/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_15/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_12/m2_390_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_14/m2_90_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_5/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_13/m2_390_n50# 018SRAM_cell1_cutPC_64x8m81_1/a_246_342#
+ 018SRAM_cell1_dummy_64x8m81_1/m2_90_n50# 018SRAM_cell1_cutPC_64x8m81_5/a_246_712#
+ VSS 018SRAM_cell1_dummy_64x8m81_14/m2_390_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_8/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_15/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_16/m2_390_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_6/m2_90_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_15/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_10/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_20/m2_90_n50#
+ 018SRAM_cell1_dummy_64x8m81_17/m2_390_n50# 018SRAM_cell1_cutPC_64x8m81_2/a_246_342#
+ 018SRAM_cell1_dummy_64x8m81_2/m2_90_n50# 018SRAM_cell1_cutPC_64x8m81_4/a_246_712#
+ 018SRAM_cell1_dummy_64x8m81_18/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_30/m2_90_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_9/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_19/m2_390_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_7/m2_90_n50# 018SRAM_cell1_dummy_64x8m81_11/m2_90_n50#
+ 018SRAM_cell1_64x8m81_0/w_n68_622# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_0/m2_390_n50#
+ 018SRAM_cell1_dummy_64x8m81_21/m2_90_n50# 018SRAM_cell1_cutPC_64x8m81_3/a_246_342#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_1/m2_390_n50# 018SRAM_cell1_dummy_64x8m81_3/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_64x8m81_31/m2_90_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_cutPC_64x8m81_0/m3_n36_330#
X018SRAM_cell1_dummy_64x8m81_30 VSUBS 018SRAM_cell1_dummy_64x8m81_30/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_30/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_31 VSUBS 018SRAM_cell1_dummy_64x8m81_31/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_31/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_20 VSUBS 018SRAM_cell1_dummy_64x8m81_20/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_20/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_22 VSUBS 018SRAM_cell1_dummy_64x8m81_22/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_22/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_21 VSUBS 018SRAM_cell1_dummy_64x8m81_21/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_21/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_11 VSUBS 018SRAM_cell1_dummy_64x8m81_11/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_11/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_10 VSUBS 018SRAM_cell1_dummy_64x8m81_10/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_10/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_23 VSUBS 018SRAM_cell1_dummy_64x8m81_23/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_23/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_12 VSUBS 018SRAM_cell1_dummy_64x8m81_12/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_12/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_24 VSUBS 018SRAM_cell1_dummy_64x8m81_24/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_24/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_13 VSUBS 018SRAM_cell1_dummy_64x8m81_13/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_13/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_25 VSUBS 018SRAM_cell1_dummy_64x8m81_25/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_25/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_14 VSUBS 018SRAM_cell1_dummy_64x8m81_14/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_14/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_26 VSUBS 018SRAM_cell1_dummy_64x8m81_26/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_26/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_15 VSUBS 018SRAM_cell1_dummy_64x8m81_15/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_15/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_cutPC_64x8m81_0 VSUBS 018SRAM_cell1_64x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_64x8m81_0/a_246_342#
+ 018SRAM_cell1_cutPC_64x8m81_7/a_246_712# 018SRAM_cell1_cutPC_64x8m81_0/m3_n36_330#
+ 018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_64x8m81_7/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_64x8m81
X018SRAM_cell1_dummy_64x8m81_27 VSUBS 018SRAM_cell1_dummy_64x8m81_27/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_27/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_16 VSUBS 018SRAM_cell1_dummy_64x8m81_16/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_16/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_0 VSUBS 018SRAM_cell1_dummy_64x8m81_0/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_0/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
Xnew_dummyrow_unit_64x8m81_0 new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_12/m2_90_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_4/m2_90_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_13/m2_90_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_5/m2_90_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_14/m2_90_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_6/m2_90_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_15/m2_90_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_7/m2_90_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_8/m2_90_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_9/m2_90_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_0/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_2/m2_390_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_1/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_3/m2_390_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_4/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_5/m2_390_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_6/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_7/m2_390_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_8/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_10/m2_390_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_9/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_0/m2_90_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_11/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_13/m2_390_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_12/m2_390_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_14/m2_390_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_1/m2_90_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_15/m2_390_n50# VSUBS new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_10/m2_90_n50#
+ new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_2/m2_90_n50# new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_11/m2_90_n50#
+ VSUBS new_dummyrow_unit_64x8m81_0/018SRAM_cell1_dummy_64x8m81_3/m2_90_n50# 018SRAM_cell1_64x8m81_1/w_n68_622#
+ new_dummyrow_unit_64x8m81
X018SRAM_cell1_cutPC_64x8m81_1 VSUBS 018SRAM_cell1_64x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_64x8m81_1/a_246_342#
+ 018SRAM_cell1_cutPC_64x8m81_5/a_246_712# 018SRAM_cell1_cutPC_64x8m81_1/m3_n36_330#
+ 018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_64x8m81_5/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_64x8m81
X018SRAM_cell1_dummy_64x8m81_28 VSUBS 018SRAM_cell1_dummy_64x8m81_28/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_28/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_17 VSUBS 018SRAM_cell1_dummy_64x8m81_17/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_17/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_1 VSUBS 018SRAM_cell1_dummy_64x8m81_1/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_1/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_cutPC_64x8m81_2 VSUBS 018SRAM_cell1_64x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_64x8m81_2/a_246_342#
+ 018SRAM_cell1_cutPC_64x8m81_4/a_246_712# 018SRAM_cell1_cutPC_64x8m81_2/m3_n36_330#
+ 018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_64x8m81_4/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_64x8m81
X018SRAM_cell1_dummy_64x8m81_29 VSUBS 018SRAM_cell1_dummy_64x8m81_29/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_29/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_18 VSUBS 018SRAM_cell1_dummy_64x8m81_18/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_18/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_2 VSUBS 018SRAM_cell1_dummy_64x8m81_2/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_2/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_cutPC_64x8m81_3 VSUBS 018SRAM_cell1_64x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_64x8m81_3/a_246_342#
+ 018SRAM_cell1_64x8m81_1/w_n68_622# 018SRAM_cell1_cutPC_64x8m81_3/m3_n36_330# 018SRAM_cell1_64x8m81_1/a_36_n42#
+ 018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_cutPC_64x8m81
X018SRAM_cell1_dummy_64x8m81_19 VSUBS 018SRAM_cell1_dummy_64x8m81_19/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_19/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_3 VSUBS 018SRAM_cell1_dummy_64x8m81_3/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_3/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_64x8m81_0 VSUBS 018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_64x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ x018SRAM_cell1_64x8m81
X018SRAM_cell1_cutPC_64x8m81_4 VSUBS 018SRAM_cell1_64x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_64x8m81_4/a_246_342#
+ 018SRAM_cell1_cutPC_64x8m81_4/a_246_712# 018SRAM_cell1_cutPC_64x8m81_4/m3_n36_330#
+ 018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_64x8m81_4/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_64x8m81
X018SRAM_cell1_dummy_64x8m81_5 VSUBS 018SRAM_cell1_dummy_64x8m81_5/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_5/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_4 VSUBS 018SRAM_cell1_dummy_64x8m81_4/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_4/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_64x8m81_1 VSUBS 018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_64x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS
+ x018SRAM_cell1_64x8m81
X018SRAM_cell1_cutPC_64x8m81_6 VSUBS 018SRAM_cell1_64x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_64x8m81_6/a_246_342#
+ 018SRAM_cell1_64x8m81_0/w_n68_622# 018SRAM_cell1_cutPC_64x8m81_6/m3_n36_330# 018SRAM_cell1_64x8m81_1/a_36_n42#
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_cutPC_64x8m81
X018SRAM_cell1_cutPC_64x8m81_5 VSUBS 018SRAM_cell1_64x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_64x8m81_5/a_246_342#
+ 018SRAM_cell1_cutPC_64x8m81_5/a_246_712# 018SRAM_cell1_cutPC_64x8m81_5/m3_n36_330#
+ 018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_64x8m81_5/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_64x8m81
X018SRAM_cell1_dummy_64x8m81_6 VSUBS 018SRAM_cell1_dummy_64x8m81_6/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_6/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_cutPC_64x8m81_7 VSUBS 018SRAM_cell1_64x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_64x8m81_7/a_246_342#
+ 018SRAM_cell1_cutPC_64x8m81_7/a_246_712# 018SRAM_cell1_cutPC_64x8m81_7/m3_n36_330#
+ 018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_64x8m81_7/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_64x8m81
X018SRAM_cell1_dummy_64x8m81_7 VSUBS 018SRAM_cell1_dummy_64x8m81_7/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_7/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_8 VSUBS 018SRAM_cell1_dummy_64x8m81_8/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_8/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
X018SRAM_cell1_dummy_64x8m81_9 VSUBS 018SRAM_cell1_dummy_64x8m81_9/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_64x8m81_9/m2_390_n50# 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_64x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_64x8m81
Xnew_dummyrow_unit_01_64x8m81_0 new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_12/m2_90_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_4/m2_90_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_13/m2_90_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_5/m2_90_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_14/m2_90_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_6/m2_90_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_15/m2_90_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_7/m2_90_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_8/m2_90_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_0/m2_390_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_9/m2_90_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_2/m2_390_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_1/m2_390_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_3/m2_390_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_5/m2_390_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_4/m2_390_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_6/m2_390_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_7/m2_390_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_0/m2_90_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_8/m2_390_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_9/m2_390_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_10/m2_390_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_11/m2_390_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_13/m2_390_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_12/m2_390_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_14/m2_390_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_1/m2_90_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_15/m2_390_n50# VSUBS
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_10/m2_90_n50# new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_2/m2_90_n50#
+ new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_11/m2_90_n50# VSUBS new_dummyrow_unit_01_64x8m81_0/018SRAM_cell1_dummy_64x8m81_3/m2_90_n50#
+ 018SRAM_cell1_64x8m81_1/w_n68_622# new_dummyrow_unit_01_64x8m81
.ends

.subckt col_64a_64x8m81_0 018SRAM_cell1_2x_64x8m81_0/018SRAM_cell1_64x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_64x8m81_97/018SRAM_cell1_64x8m81_1/a_444_n42# 018SRAM_cell1_2x_64x8m81_45/018SRAM_cell1_64x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_64x8m81_46/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_88/018SRAM_cell1_64x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_64x8m81_94/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_7/018SRAM_cell1_64x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_64x8m81_7/018SRAM_cell1_64x8m81_1/a_444_n42# 018SRAM_cell1_2x_64x8m81_90/018SRAM_cell1_64x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_64x8m81_6/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_64x8m81_5/018SRAM_cell1_64x8m81_1/a_444_n42# 018SRAM_cell1_2x_64x8m81_32/018SRAM_cell1_64x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_64x8m81_36/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_87/018SRAM_cell1_64x8m81_1/a_444_n42# 018SRAM_cell1_2x_64x8m81_45/018SRAM_cell1_64x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_64x8m81_93/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_35/018SRAM_cell1_64x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_64x8m81_92/018SRAM_cell1_64x8m81_1/a_444_n42# 018SRAM_cell1_2x_64x8m81_96/018SRAM_cell1_64x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_64x8m81_57/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_57/018SRAM_cell1_64x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_64x8m81_92/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_34/018SRAM_cell1_64x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_64x8m81_2/018SRAM_cell1_64x8m81_1/a_444_n42# 018SRAM_cell1_2x_64x8m81_56/018SRAM_cell1_64x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_64x8m81_3/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_46/018SRAM_cell1_64x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_64x8m81_1/018SRAM_cell1_64x8m81_1/a_444_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_88/018SRAM_cell1_64x8m81_1/a_444_n42# 018SRAM_cell1_2x_64x8m81_34/018SRAM_cell1_64x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_64x8m81_89/018SRAM_cell1_64x8m81_1/a_444_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_91/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_8/018SRAM_cell1_64x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_64x8m81_2/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_98/018SRAM_cell1_64x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_4/018SRAM_cell1_64x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_64x8m81_47/018SRAM_cell1_64x8m81_1/a_444_n42# 018SRAM_cell1_2x_64x8m81_6/018SRAM_cell1_64x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# 018SRAM_cell1_2x_64x8m81_90/018SRAM_cell1_64x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_64x8m81_96/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_64x8m81_32/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_1/018SRAM_cell1_64x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_64x8m81_93/018SRAM_cell1_64x8m81_1/a_444_n42# 018SRAM_cell1_2x_64x8m81_98/018SRAM_cell1_64x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_64x8m81_5/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_94/018SRAM_cell1_64x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_444_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_35/018SRAM_cell1_64x8m81_1/a_444_n42# 018SRAM_cell1_2x_64x8m81_3/018SRAM_cell1_64x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# 018SRAM_cell1_2x_64x8m81_36/018SRAM_cell1_64x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_64x8m81_8/018SRAM_cell1_64x8m81_1/a_444_n42# 018SRAM_cell1_2x_64x8m81_33/018SRAM_cell1_64x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_64x8m81_89/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_91/018SRAM_cell1_64x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_87/018SRAM_cell1_64x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_64x8m81_47/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_0/018SRAM_cell1_64x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_64x8m81_97/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_56/018SRAM_cell1_64x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_4/018SRAM_cell1_64x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_64x8m81_33/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
X018SRAM_cell1_2x_64x8m81_1 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_1/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_1/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_2 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_2/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_2/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_3 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_3/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_3/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_4 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_4/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_4/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_5 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_5/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_5/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_6 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_6/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_6/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_7 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_7/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_7/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_8 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_8/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_8/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_9 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_90 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_90/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_90/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_80 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_88/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_88/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_91 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_91/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_91/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_70 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_5/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_5/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_81 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_89/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_89/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_92 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_92/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_92/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_120 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_46/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_46/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_60 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_5/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_5/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_82 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_90/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_90/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_71 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_1/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_1/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_93 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_93/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_93/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_110 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_0/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_0/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_121 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_47/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_47/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_61 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_4/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_4/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_50 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_7/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_7/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_83 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_91/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_91/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_72 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_2/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_2/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_94 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_94/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_94/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_111 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_6/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_6/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_100 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_56/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_56/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_122 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_32/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_32/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_62 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_3/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_3/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_51 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_6/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_6/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_40 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_90/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_90/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_95 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_8/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_8/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_84 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_92/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_92/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_73 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_3/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_3/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_112 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_46/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_46/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_101 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_57/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_57/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_123 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_33/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_33/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_63 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_1/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_1/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_52 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_96/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_96/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_41 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_91/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_91/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_85 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_93/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_93/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_30 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_94/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_94/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_96 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_96/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_96/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_74 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_4/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_4/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_113 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_47/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_47/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_102 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_0/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_0/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_124 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_34/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_34/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_20 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_34/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_34/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_53 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_97/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_97/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_42 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_92/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_92/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_64 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_7/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_7/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_86 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_94/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_94/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_31 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_87/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_87/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_97 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_97/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_97/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_75 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_5/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_5/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_114 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_32/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_32/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_103 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_6/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_6/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_125 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_35/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_35/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_54 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_98/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_98/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_43 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_93/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_93/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_32 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_32/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_32/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_65 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_21 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_35/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_35/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_10 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_96/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_96/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_98 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_98/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_98/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_76 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_7/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_7/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_87 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_87/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_87/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_115 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_33/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_33/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_126 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_36/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_36/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_104 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_96/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_96/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_55 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_44 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_94/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_94/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_33 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_33/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_33/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_66 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_1/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_1/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_22 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_36/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_36/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_11 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_97/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_97/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_99 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_77 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_8/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_8/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_88 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_88/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_88/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_116 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_34/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_34/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_127 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_45/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_45/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_105 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_97/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_97/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_56 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_56/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_56/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_45 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_45/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_45/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_34 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_34/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_34/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_67 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_2/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_2/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_23 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_45/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_45/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_12 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_98/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_98/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_78 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_89 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_89/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_89/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_106 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_98/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_98/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_117 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_35/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_35/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_57 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_57/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_57/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_35 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_35/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_35/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_46 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_46/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_46/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_68 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_3/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_3/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_79 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_87/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_87/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_24 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_88/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_88/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_13 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_118 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_36/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_36/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_107 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_58 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_0/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_0/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_36 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_36/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_36/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_47 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_47/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_47/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_69 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_4/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_4/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_25 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_89/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_89/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_14 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_56/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_56/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_108 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_56/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_56/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_119 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_45/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_45/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_99/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_59 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_2/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_2/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_48 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_37 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_87/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_87/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_26 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_90/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_90/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_15 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_57/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_57/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_109 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_57/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_57/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_95/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_49 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_8/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_8/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_38 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_88/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_88/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_16 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_46/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_46/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_27 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_91/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_91/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_39 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_89/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_89/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_63/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_17 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_47/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_47/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_28 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_92/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_92/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_18 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_32/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_32/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_29 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_93/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_93/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_19 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_33/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_33/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
X018SRAM_cell1_2x_64x8m81_0 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_0/018SRAM_cell1_64x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_0/018SRAM_cell1_64x8m81_1/a_36_n42# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/a_n36_52# 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_64x8m81_9/018SRAM_cell1_64x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_2x_64x8m81
.ends

.subckt lcol4_64_64x8m81 pcb[2] pcb[3] pcb[0] pcb[1] vdd WEN[3] WEN[2] WEN[1] WEN[0]
+ WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] ypass[0] ypass[1] ypass[2] ypass[3]
+ ypass[4] ypass[5] GWEN din[0] din[1] din[2] q[1] b[1] b[4] b[7] b[10] b[13] b[16]
+ b[19] b[22] b[25] b[28] b[31] din[3] q[0] q[2] q[3] b[29] b[26] b[23] b[20] b[17]
+ b[14] b[11] b[8] b[5] b[2] bb[0] bb[1] bb[2] bb[3] bb[4] bb[5] bb[6] bb[7] bb[8]
+ bb[9] bb[10] bb[11] bb[12] bb[13] bb[14] bb[15] bb[16] bb[17] bb[18] bb[19] bb[20]
+ bb[21] bb[22] bb[23] bb[24] bb[25] bb[26] bb[27] bb[28] bb[29] bb[30] bb[31] b[30]
+ b[27] b[24] b[15] b[12] b[9] b[21] b[0] b[3] b[6] b[18] a_15488_27175# a_15488_27950#
+ ldummy_64x4_64x8m81_0/VSS saout_R_m2_64x8m81_0/wen_wm1_64x8m81_0/wen a_4688_27175#
+ a_15248_27175# a_4688_27950# men a_15248_27950# a_4448_27175# saout_m2_64x8m81_1/mux821_64x8m81_0/a_656_7735#
+ ypass[6] a_4448_27950# ypass[7] saout_R_m2_64x8m81_1/sa_64x8m81_0/pcb saout_m2_64x8m81_1/sa_64x8m81_0/pcb
+ saout_R_m2_64x8m81_0/sa_64x8m81_0/pcb saout_m2_64x8m81_0/pcb GWE saout_m2_64x8m81_0/WEN
+ VSS VDD
Xdcap_103_novia_64x8m81_0[0] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[1] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[2] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[3] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[4] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[5] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[6] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[7] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[8] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[9] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[10] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[11] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[12] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[13] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[14] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[15] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[16] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[17] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[18] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[19] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[20] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[21] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[22] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[23] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[24] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[25] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[26] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[27] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[28] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[29] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[30] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[31] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[32] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[33] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[34] VDD VDD VSS dcap_103_novia_64x8m81
Xdcap_103_novia_64x8m81_0[35] VDD VDD VSS dcap_103_novia_64x8m81
Xsaout_R_m2_64x8m81_0 saout_R_m2_64x8m81_0/pcb saout_R_m2_64x8m81_0/datain saout_R_m2_64x8m81_0/WEN
+ ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7] men ypass[0] GWEN
+ b[0] saout_R_m2_64x8m81_0/q bb[1] saout_R_m2_64x8m81_0/sa_64x8m81_0/wep VSS GWE
+ bb[2] b[3] bb[5] ypass[7] bb[0] VSS saout_m2_64x8m81_1/mux821_64x8m81_0/a_656_7735#
+ b[7] GWEN a_15714_27175# a_15488_27175# b[2] b[6] bb[3] a_15714_27950# a_15488_27950#
+ b[5] b[1] bb[4] men b[4] ypass[0] bb[6] ypass[2] ypass[1] saout_R_m2_64x8m81_0/wen_wm1_64x8m81_0/wen
+ ypass[5] VDD bb[7] ypass[6] saout_R_m2_64x8m81_0/sa_64x8m81_0/pcb saout_R_m2_64x8m81_0/sacntl_2_64x8m81_0/a_4718_983#
+ b[5] ypass[3] ypass[4] VSS VDD VDD VDD saout_R_m2_64x8m81
Xsaout_R_m2_64x8m81_1 saout_R_m2_64x8m81_1/pcb saout_R_m2_64x8m81_1/datain saout_R_m2_64x8m81_1/WEN
+ ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7] men ypass[0] GWEN
+ b[16] saout_R_m2_64x8m81_1/q bb[17] saout_R_m2_64x8m81_1/sa_64x8m81_0/wep VSS GWE
+ bb[18] b[19] bb[21] ypass[7] bb[16] VSS saout_m2_64x8m81_1/mux821_64x8m81_0/a_656_7735#
+ b[23] GWEN a_4914_27175# a_4688_27175# b[18] b[22] bb[19] a_4914_27950# a_4688_27950#
+ b[21] b[17] bb[20] men b[20] ypass[0] bb[22] ypass[2] ypass[1] saout_R_m2_64x8m81_1/wen_wm1_64x8m81_0/wen
+ ypass[5] VDD bb[23] ypass[6] saout_R_m2_64x8m81_1/sa_64x8m81_0/pcb VSS saout_R_m2_64x8m81_1/mux821_64x8m81_0/ypass_gate_64x8m81_4/b
+ ypass[3] ypass[4] VSS VDD VDD VDD saout_R_m2_64x8m81
Xsaout_m2_64x8m81_0 saout_m2_64x8m81_0/pcb saout_m2_64x8m81_0/datain saout_m2_64x8m81_0/WEN
+ ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7] men ypass[0] GWEN
+ bb[29] bb[30] b[24] saout_m2_64x8m81_0/q a_4223_27175# a_4448_27175# saout_m2_64x8m81_0/sa_64x8m81_0/wep
+ a_4223_27950# a_4448_27950# VSS GWE saout_m2_64x8m81_0/mux821_64x8m81_0/a_4992_424#
+ b[28] bb[26] bb[31] VSS saout_m2_64x8m81_1/mux821_64x8m81_0/a_656_7735# GWEN ypass[7]
+ b[31] b[29] b[25] bb[28] b[26] b[30] bb[27] b[27] saout_m2_64x8m81_0/mux821_64x8m81_0/ypass_gate_a_64x8m81_0/a_n80_n10#
+ ypass[0] bb[25] ypass[2] ypass[1] VDD bb[24] saout_m2_64x8m81_0/pcb saout_m2_64x8m81_0/sacntl_2_64x8m81_0/a_4718_983#
+ men ypass[5] VDD ypass[3] ypass[4] saout_m2_64x8m81_0/mux821_64x8m81_0/ypass_gate_a_64x8m81_0/b
+ ypass[6] VSS VDD VDD saout_m2_64x8m81
Xldummy_64x4_64x8m81_0 b[5] WL[3] b[3] bb[25] bb[13] WL[5] bb[2] b[16] bb[22] VSS
+ bb[3] WL[7] b[1] bb[20] WL[6] b[6] bb[0] b[21] WL[4] bb[8] b[12] b[19] b[26] WL[0]
+ b[9] bb[18] b[24] VSS WL[2] VDD bb[10] b[2] b[17] b[4] bb[16] b[14] bb[24] b[25]
+ bb[25] VSS b[27] VDD bb[26] bb[1] b[29] bb[5] bb[28] bb[11] b[22] b[31] bb[30] bb[15]
+ b[26] b[23] b[31] VSS VDD b[11] b[0] b[23] b[13] bb[3] bb[13] bb[12] b[20] b[22]
+ bb[27] bb[14] bb[27] b[15] b[8] b[7] b[2] bb[29] b[12] bb[21] b[20] bb[29] b[7]
+ bb[18] bb[9] b[17] bb[6] bb[1] bb[16] bb[4] b[14] b[28] bb[24] bb[19] b[5] bb[21]
+ b[25] b[28] b[3] bb[2] bb[26] b[0] b[1] b[27] bb[15] bb[0] bb[19] b[29] b[18] b[30]
+ bb[28] b[30] bb[8] VSS VDD bb[7] bb[10] b[9] bb[30] b[8] b[11] bb[7] b[13] bb[31]
+ bb[17] bb[12] VSS b[6] VDD ldummy_64x4_64x8m81_0/VSS bb[14] bb[9] b[15] bb[22] b[16]
+ bb[23] b[10] b[18] bb[20] VSS b[4] VDD b[21] bb[31] b[10] b[19] b[24] bb[11] VDD
+ bb[6] bb[17] VSS bb[4] bb[5] VSS bb[23] VDD WL[1] ldummy_64x4_64x8m81
Xsaout_m2_64x8m81_1 saout_m2_64x8m81_1/pcb saout_m2_64x8m81_1/datain saout_m2_64x8m81_1/WEN
+ ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7] men ypass[0] GWEN
+ bb[13] bb[14] b[8] saout_m2_64x8m81_1/q a_15023_27175# a_15248_27175# saout_m2_64x8m81_1/sa_64x8m81_0/wep
+ a_15023_27950# a_15248_27950# VSS GWE VSS b[12] bb[10] bb[15] VSS saout_m2_64x8m81_1/mux821_64x8m81_0/a_656_7735#
+ GWEN ypass[7] b[15] b[13] b[9] bb[12] b[10] b[14] bb[11] b[11] VSS ypass[0] bb[9]
+ ypass[2] ypass[1] VDD bb[8] saout_m2_64x8m81_1/sa_64x8m81_0/pcb VSS men ypass[5]
+ VDD ypass[3] ypass[4] saout_m2_64x8m81_1/mux821_64x8m81_0/ypass_gate_a_64x8m81_0/b
+ ypass[6] VSS VDD VDD saout_m2_64x8m81
Xcol_64a_64x8m81_0_0 bb[9] b[14] bb[24] b[31] bb[17] bb[23] bb[7] b[7] b[19] bb[8]
+ b[12] b[1] bb[29] b[25] WL[3] bb[16] b[24] b[22] bb[26] b[21] bb[15] bb[10] b[10]
+ bb[21] b[27] bb[0] b[11] bb[3] bb[31] bb[4] WL[6] b[17] bb[27] bb[18] WL[1] b[20]
+ b[6] b[0] bb[13] bb[12] b[2] b[30] b[8] WL[4] bb[19] b[15] bb[5] b[29] b[4] bb[22]
+ b[13] bb[1] b[23] b[5] WL[0] b[26] b[3] WL[2] bb[25] bb[6] bb[28] b[18] bb[20] WL[7]
+ b[16] bb[30] b[9] bb[14] bb[11] WL[5] bb[2] b[28] VSS VDD col_64a_64x8m81_0
.ends

.subckt gf180mcu_fd_ip_sram__sram64x8m8wm1 VSS CLK D[0] A[2] A[1] A[0] Q[2] Q[3] CEN
+ A[5] A[4] WEN[3] D[7] Q[7] D[3] D[1] D[2] A[3] Q[1] Q[6] D[5] Q[4] WEN[5] WEN[2]
+ WEN[1] WEN[4] WEN[7] WEN[6] D[4] D[6] Q[5] Q[0] GWEN WEN[0]
Xcontrol_512x8_64x8m81_0 rcol4_64_64x8m81_0/GWE GWEN VSS VSS rcol4_64_64x8m81_0/ypass[7]
+ rcol4_64_64x8m81_0/ypass[6] rcol4_64_64x8m81_0/ypass[5] rcol4_64_64x8m81_0/ypass[4]
+ rcol4_64_64x8m81_0/ypass[3] rcol4_64_64x8m81_0/ypass[1] rcol4_64_64x8m81_0/ypass[0]
+ lcol4_64_64x8m81_0/ypass[0] lcol4_64_64x8m81_0/ypass[1] lcol4_64_64x8m81_0/ypass[2]
+ lcol4_64_64x8m81_0/ypass[3] lcol4_64_64x8m81_0/ypass[6] lcol4_64_64x8m81_0/ypass[5]
+ lcol4_64_64x8m81_0/ypass[4] lcol4_64_64x8m81_0/ypass[7] rcol4_64_64x8m81_0/tblhl
+ control_512x8_64x8m81_0/xb[3] control_512x8_64x8m81_0/xb[2] control_512x8_64x8m81_0/xb[0]
+ xdec8_64_64x8m81_0/xa[7] xdec8_64_64x8m81_0/xa[5] xdec8_64_64x8m81_0/xa[4] xdec8_64_64x8m81_0/xa[3]
+ xdec8_64_64x8m81_0/xa[2] A[0] control_512x8_64x8m81_0/xb[1] control_512x8_64x8m81_0/xc[3]
+ control_512x8_64x8m81_0/xc[1] control_512x8_64x8m81_0/xc[2] control_512x8_64x8m81_0/xc[0]
+ xdec8_64_64x8m81_0/xa[0] xdec8_64_64x8m81_0/xa[1] VSS VSS CLK A[2] A[1] VSS A[3]
+ A[4] A[5] VSS lcol4_64_64x8m81_0/ypass[2] rcol4_64_64x8m81_0/tblhl rcol4_64_64x8m81_0/GWEN
+ control_512x8_64x8m81_0/gen_512x8_64x8m81_0/wen_v2_64x8m81_0/nmos_5p0431058998329_64x8m81_4/D
+ CEN xdec8_64_64x8m81_0/xa[6] rcol4_64_64x8m81_0/ypass[2] VSS xdec8_64_64x8m81_0/men
+ VSS VSS VSS control_512x8_64x8m81
Xrcol4_64_64x8m81_0 rcol4_64_64x8m81_0/pcb[6] rcol4_64_64x8m81_0/pcb[7] rcol4_64_64x8m81_0/pcb[4]
+ VSS WEN[7] WEN[4] rcol4_64_64x8m81_0/pcb[5] WEN[6] WEN[5] rcol4_64_64x8m81_0/WL[6]
+ rcol4_64_64x8m81_0/WL[5] rcol4_64_64x8m81_0/ypass[1] rcol4_64_64x8m81_0/ypass[2]
+ rcol4_64_64x8m81_0/ypass[3] rcol4_64_64x8m81_0/ypass[4] rcol4_64_64x8m81_0/ypass[5]
+ rcol4_64_64x8m81_0/ypass[6] rcol4_64_64x8m81_0/DWL rcol4_64_64x8m81_0/tblhl rcol4_64_64x8m81_0/GWEN
+ rcol4_64_64x8m81_0/ypass[0] rcol4_64_64x8m81_0/WL[0] rcol4_64_64x8m81_0/WL[2] rcol4_64_64x8m81_0/WL[3]
+ rcol4_64_64x8m81_0/WL[4] rcol4_64_64x8m81_0/WL[7] rcol4_64_64x8m81_0/WL[1] rcol4_64_64x8m81_0/ypass[7]
+ D[4] D[7] Q[5] Q[6] Q[7] D[5] D[6] Q[4] VSS xdec8_64_64x8m81_0/men rcol4_64_64x8m81_0/WL[0]
+ rcol4_64_64x8m81_0/saout_R_m2_64x8m81_1/pcb VSS rcol4_64_64x8m81_0/WL[1] rcol4_64_64x8m81_0/WL[2]
+ rcol4_64_64x8m81_0/WL[3] rcol4_64_64x8m81_0/WL[4] rcol4_64_64x8m81_0/WL[5] rcol4_64_64x8m81_0/WL[6]
+ rcol4_64_64x8m81_0/WL[7] VSS rcol4_64_64x8m81_0/DWL VSS VSS VSS WEN[7] VSS VSS VSS
+ VSS VSS VSS VSS rcol4_64_64x8m81_0/saout_R_m2_64x8m81_1/pcb rcol4_64_64x8m81_0/saout_m2_64x8m81_1/sa_64x8m81_0/pcb
+ rcol4_64_64x8m81_0/saout_R_m2_64x8m81_0/sa_64x8m81_0/pcb rcol4_64_64x8m81_0/saout_m2_64x8m81_0/pcb
+ rcol4_64_64x8m81_0/GWE VSS VSS rcol4_64_64x8m81
Xxdec8_64_64x8m81_0 rcol4_64_64x8m81_0/DWL rcol4_64_64x8m81_0/WL[6] rcol4_64_64x8m81_0/WL[1]
+ lcol4_64_64x8m81_0/WL[6] lcol4_64_64x8m81_0/WL[7] lcol4_64_64x8m81_0/WL[2] lcol4_64_64x8m81_0/WL[3]
+ lcol4_64_64x8m81_0/WL[4] lcol4_64_64x8m81_0/WL[5] lcol4_64_64x8m81_0/WL[0] xdec8_64_64x8m81_0/DLWL
+ xdec8_64_64x8m81_0/xa[7] xdec8_64_64x8m81_0/xa[6] xdec8_64_64x8m81_0/xa[5] xdec8_64_64x8m81_0/xa[4]
+ xdec8_64_64x8m81_0/xa[0] xdec8_64_64x8m81_0/xa[3] xdec8_64_64x8m81_0/xa[2] xdec8_64_64x8m81_0/xa[1]
+ rcol4_64_64x8m81_0/WL[4] rcol4_64_64x8m81_0/WL[2] rcol4_64_64x8m81_0/WL[0] xdec8_64_64x8m81_0/men
+ lcol4_64_64x8m81_0/WL[1] rcol4_64_64x8m81_0/WL[7] rcol4_64_64x8m81_0/WL[5] rcol4_64_64x8m81_0/WL[3]
+ VSS VSS xdec8_64_64x8m81
Xlcol4_64_64x8m81_0 lcol4_64_64x8m81_0/pcb[2] lcol4_64_64x8m81_0/pcb[3] lcol4_64_64x8m81_0/pcb[0]
+ lcol4_64_64x8m81_0/pcb[1] VSS WEN[0] WEN[1] WEN[2] WEN[3] lcol4_64_64x8m81_0/WL[7]
+ lcol4_64_64x8m81_0/WL[6] lcol4_64_64x8m81_0/WL[5] lcol4_64_64x8m81_0/WL[4] lcol4_64_64x8m81_0/WL[3]
+ lcol4_64_64x8m81_0/WL[2] lcol4_64_64x8m81_0/WL[1] lcol4_64_64x8m81_0/WL[0] lcol4_64_64x8m81_0/ypass[0]
+ lcol4_64_64x8m81_0/ypass[1] lcol4_64_64x8m81_0/ypass[2] lcol4_64_64x8m81_0/ypass[3]
+ lcol4_64_64x8m81_0/ypass[4] lcol4_64_64x8m81_0/ypass[5] rcol4_64_64x8m81_0/GWEN
+ D[0] D[1] D[2] Q[1] lcol4_64_64x8m81_0/b[1] lcol4_64_64x8m81_0/b[4] lcol4_64_64x8m81_0/b[7]
+ lcol4_64_64x8m81_0/b[10] lcol4_64_64x8m81_0/b[13] lcol4_64_64x8m81_0/b[16] lcol4_64_64x8m81_0/b[19]
+ lcol4_64_64x8m81_0/b[22] lcol4_64_64x8m81_0/b[25] lcol4_64_64x8m81_0/b[28] lcol4_64_64x8m81_0/b[31]
+ D[3] Q[0] Q[2] Q[3] lcol4_64_64x8m81_0/b[29] lcol4_64_64x8m81_0/b[26] lcol4_64_64x8m81_0/b[23]
+ lcol4_64_64x8m81_0/b[20] lcol4_64_64x8m81_0/b[17] lcol4_64_64x8m81_0/b[14] lcol4_64_64x8m81_0/b[11]
+ lcol4_64_64x8m81_0/b[8] lcol4_64_64x8m81_0/b[5] lcol4_64_64x8m81_0/b[2] lcol4_64_64x8m81_0/bb[0]
+ lcol4_64_64x8m81_0/bb[1] lcol4_64_64x8m81_0/bb[2] lcol4_64_64x8m81_0/bb[3] lcol4_64_64x8m81_0/bb[4]
+ lcol4_64_64x8m81_0/bb[5] lcol4_64_64x8m81_0/bb[6] lcol4_64_64x8m81_0/bb[7] lcol4_64_64x8m81_0/bb[8]
+ lcol4_64_64x8m81_0/bb[9] lcol4_64_64x8m81_0/bb[10] lcol4_64_64x8m81_0/bb[11] lcol4_64_64x8m81_0/bb[12]
+ lcol4_64_64x8m81_0/bb[13] lcol4_64_64x8m81_0/bb[14] lcol4_64_64x8m81_0/bb[15] lcol4_64_64x8m81_0/bb[16]
+ lcol4_64_64x8m81_0/bb[17] lcol4_64_64x8m81_0/bb[18] lcol4_64_64x8m81_0/bb[19] lcol4_64_64x8m81_0/bb[20]
+ lcol4_64_64x8m81_0/bb[21] lcol4_64_64x8m81_0/bb[22] lcol4_64_64x8m81_0/bb[23] lcol4_64_64x8m81_0/bb[24]
+ lcol4_64_64x8m81_0/bb[25] lcol4_64_64x8m81_0/bb[26] lcol4_64_64x8m81_0/bb[27] lcol4_64_64x8m81_0/bb[28]
+ lcol4_64_64x8m81_0/bb[29] lcol4_64_64x8m81_0/bb[30] lcol4_64_64x8m81_0/bb[31] lcol4_64_64x8m81_0/b[30]
+ lcol4_64_64x8m81_0/b[27] lcol4_64_64x8m81_0/b[24] lcol4_64_64x8m81_0/b[15] lcol4_64_64x8m81_0/b[12]
+ lcol4_64_64x8m81_0/b[9] lcol4_64_64x8m81_0/b[21] lcol4_64_64x8m81_0/b[0] lcol4_64_64x8m81_0/b[3]
+ lcol4_64_64x8m81_0/b[6] lcol4_64_64x8m81_0/b[18] VSS VSS VSS WEN[3] VSS VSS VSS
+ xdec8_64_64x8m81_0/men VSS VSS VSS lcol4_64_64x8m81_0/ypass[6] VSS lcol4_64_64x8m81_0/ypass[7]
+ lcol4_64_64x8m81_0/saout_R_m2_64x8m81_1/sa_64x8m81_0/pcb lcol4_64_64x8m81_0/saout_m2_64x8m81_1/sa_64x8m81_0/pcb
+ lcol4_64_64x8m81_0/saout_R_m2_64x8m81_0/sa_64x8m81_0/pcb lcol4_64_64x8m81_0/saout_m2_64x8m81_0/pcb
+ rcol4_64_64x8m81_0/GWE WEN[0] VSS VSS lcol4_64_64x8m81
.ends

