// //#############################################################################
// //# Function: Positive edge-triggered inverting static D-type flop-flop       #
// //#           with scan input.                                                #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_sdffqn #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      si,
//     input      se,
//     input      clk,
//     output reg qn
// );
// 
//     always @(posedge clk) qn <= se ? ~si : ~d;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_sdffqn.v:11.1-23.10" *)
module la_sdffqn (
    d,
    si,
    se,
    clk,
    qn
);
  (* src = "inputs/la_sdffqn.v:21.5-21.47" *)
  wire _0_;
  wire _1_;
  (* unused_bits = "0" *)
  wire _2_;
  wire _3_;
  (* src = "inputs/la_sdffqn.v:17.16-17.19" *)
  input clk;
  wire clk;
  (* src = "inputs/la_sdffqn.v:14.16-14.17" *)
  input d;
  wire d;
  (* src = "inputs/la_sdffqn.v:18.16-18.18" *)
  output qn;
  wire qn;
  (* src = "inputs/la_sdffqn.v:16.16-16.18" *)
  input se;
  wire se;
  (* src = "inputs/la_sdffqn.v:15.16-15.18" *)
  input si;
  wire si;
  sg13g2_nand2b_1 _4_ (
      .A_N(si),
      .B  (se),
      .Y  (_1_)
  );
  sg13g2_o21ai_1 _5_ (
      .A1(d),
      .A2(se),
      .B1(_1_),
      .Y (_0_)
  );
  (* src = "inputs/la_sdffqn.v:21.5-21.47" *)
  sg13g2_dfrbp_1 _6_ (
      .CLK(clk),
      .D(_0_),
      .Q(qn),
      .Q_N(_2_),
      .RESET_B(_3_)
  );
  sg13g2_tiehi _7_ (.L_HI(_3_));
endmodule
