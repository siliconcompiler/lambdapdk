// //#############################################################################
// //# Function: 4-Input Exclusive-Nor Gate                                      #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_xnor4 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     input  b,
//     input  c,
//     input  d,
//     output z
// );
// 
//   assign z = ~(a ^ b ^ c ^ d);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_xnor4.v:10.1-22.10" *)
module la_xnor4 (
    a,
    b,
    c,
    d,
    z
);
  wire _0_;
  wire _1_;
  (* src = "inputs/la_xnor4.v:13.12-13.13" *)
  input a;
  wire a;
  (* src = "inputs/la_xnor4.v:14.12-14.13" *)
  input b;
  wire b;
  (* src = "inputs/la_xnor4.v:15.12-15.13" *)
  input c;
  wire c;
  (* src = "inputs/la_xnor4.v:16.12-16.13" *)
  input d;
  wire d;
  (* src = "inputs/la_xnor4.v:17.12-17.13" *)
  output z;
  wire z;
  XNOR2_X2 _2_ (
      .A (c),
      .B (d),
      .ZN(_0_)
  );
  XNOR2_X2 _3_ (
      .A (b),
      .B (a),
      .ZN(_1_)
  );
  XNOR2_X2 _4_ (
      .A (_0_),
      .B (_1_),
      .ZN(z)
  );
endmodule
