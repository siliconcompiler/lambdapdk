// //#############################################################################
// //# Function: And-Or (ao222) Gate                                             #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_ao222 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a0,
//     input  a1,
//     input  b0,
//     input  b1,
//     input  c0,
//     input  c1,
//     output z
// );
// 
//     assign z = (a0 & a1) | (b0 & b1) | (c0 & c1);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
module la_ao222 (
    a0,
    a1,
    b0,
    b1,
    c0,
    c1,
    z
);
  wire _0_;
  wire _1_;
  (* src = "generated" *)
  input a0;
  wire a0;
  (* src = "generated" *)
  input a1;
  wire a1;
  (* src = "generated" *)
  input b0;
  wire b0;
  (* src = "generated" *)
  input b1;
  wire b1;
  (* src = "generated" *)
  input c0;
  wire c0;
  (* src = "generated" *)
  input c1;
  wire c1;
  (* src = "generated" *)
  output z;
  wire z;
  sg13g2_nand2_1 _2_ (
      .A(b1),
      .B(b0),
      .Y(_0_)
  );
  sg13g2_a22oi_1 _3_ (
      .A1(c1),
      .A2(c0),
      .B1(a1),
      .B2(a0),
      .Y (_1_)
  );
  sg13g2_nand2_1 _4_ (
      .A(_0_),
      .B(_1_),
      .Y(z)
  );
endmodule
