// //#############################################################################
// //# Function: And-Or-Inverter (aoi21) Gate                                    #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_aoi21 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a0,
//     input  a1,
//     input  b0,
//     output z
// );
// 
//     assign z = ~((a0 & a1) | b0);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
(* keep_hierarchy *)
module la_aoi21 (
    a0,
    a1,
    b0,
    z
);
  (* src = "generated" *)
  input a0;
  wire a0;
  (* src = "generated" *)
  input a1;
  wire a1;
  (* src = "generated" *)
  input b0;
  wire b0;
  (* src = "generated" *)
  output z;
  wire z;
  gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _0_ (
      .A1(a1),
      .A2(a0),
      .B (b0),
      .ZN(z)
  );
endmodule
