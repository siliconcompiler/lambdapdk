// //#############################################################################
// //# Function: Synchronizer with async reset                                   #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// module la_drsync #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  clk,    // clock
//     input  in,     // input data
//     input  nreset, // async active low reset
//     output out     // synchronized data
// );
// 
//     localparam STAGES = 2;
// 
//     reg [STAGES-1:0] shiftreg;
// 
//     always @(posedge clk or negedge nreset)
//         if (!nreset) shiftreg[STAGES-1:0] <= 'b0;
//         else shiftreg[STAGES-1:0] <= {shiftreg[STAGES-2:0], in};
// 
//     assign out = shiftreg[STAGES-1];
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* dynports =  1  *)
(* top =  1  *)
(* src = "generated" *)
(* keep_hierarchy *)
module la_drsync (
    clk,
    in,
    nreset,
    out
);
  (* unused_bits = "0" *)
  wire _0_;
  (* unused_bits = "0" *)
  wire _1_;
  (* src = "generated" *)
  input clk;
  wire clk;
  (* src = "generated" *)
  input in;
  wire in;
  (* src = "generated" *)
  input nreset;
  wire nreset;
  (* src = "generated" *)
  output out;
  wire out;
  (* src = "generated" *)
  wire \shiftreg[0] ;
  (* src = "generated" *)
  DFFR_X1 _2_ (
      .CK(clk),
      .D (in),
      .Q (\shiftreg[0] ),
      .QN(_1_),
      .RN(nreset)
  );
  (* src = "generated" *)
  DFFR_X1 _3_ (
      .CK(clk),
      .D (\shiftreg[0] ),
      .Q (out),
      .QN(_0_),
      .RN(nreset)
  );
endmodule
