VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO ALIGNMENT
  CLASS BLOCK ;
  SYMMETRY X Y ;
  SIZE 80.000 BY 80.000 ;
  ORIGIN 40.000 40.000 ;
  OBS
    LAYER M1 ;
    POLYGON -16.568 -40.000 -40.000 -16.568 -40.000 16.568 -16.568 40.000 0.000 40.000 0.000 32.000 -13.256 32.000 -32.000 13.256 -32.000 -13.256 -13.256 -32.000 13.256 -32.000 32.000 -13.256 32.000 13.256 13.256 32.000 0.000 32.000 0.000 40.000 16.568 40.000 40.000 16.568 40.000 -16.568 16.568 -40.000 ;
    LAYER M2 ;
    POLYGON -16.568 -40.000 -40.000 -16.568 -40.000 16.568 -16.568 40.000 0.000 40.000 0.000 32.000 -13.256 32.000 -32.000 13.256 -32.000 -13.256 -13.256 -32.000 13.256 -32.000 32.000 -13.256 32.000 13.256 13.256 32.000 0.000 32.000 0.000 40.000 16.568 40.000 40.000 16.568 40.000 -16.568 16.568 -40.000 ;
    LAYER M3 ;
    POLYGON -16.568 -40.000 -40.000 -16.568 -40.000 16.568 -16.568 40.000 0.000 40.000 0.000 32.000 -13.256 32.000 -32.000 13.256 -32.000 -13.256 -13.256 -32.000 13.256 -32.000 32.000 -13.256 32.000 13.256 13.256 32.000 0.000 32.000 0.000 40.000 16.568 40.000 40.000 16.568 40.000 -16.568 16.568 -40.000 ;
    LAYER M4 ;
    POLYGON -16.568 -40.000 -40.000 -16.568 -40.000 16.568 -16.568 40.000 0.000 40.000 0.000 32.000 -13.256 32.000 -32.000 13.256 -32.000 -13.256 -13.256 -32.000 13.256 -32.000 32.000 -13.256 32.000 13.256 13.256 32.000 0.000 32.000 0.000 40.000 16.568 40.000 40.000 16.568 40.000 -16.568 16.568 -40.000 ;
    LAYER M5 ;
    POLYGON -16.568 -40.000 -40.000 -16.568 -40.000 16.568 -16.568 40.000 0.000 40.000 0.000 32.000 -13.256 32.000 -32.000 13.256 -32.000 -13.256 -13.256 -32.000 13.256 -32.000 32.000 -13.256 32.000 13.256 13.256 32.000 0.000 32.000 0.000 40.000 16.568 40.000 40.000 16.568 40.000 -16.568 16.568 -40.000 ;
    LAYER M6 ;
    POLYGON -16.568 -40.000 -40.000 -16.568 -40.000 16.568 -16.568 40.000 0.000 40.000 0.000 32.000 -13.256 32.000 -32.000 13.256 -32.000 -13.256 -13.256 -32.000 13.256 -32.000 32.000 -13.256 32.000 13.256 13.256 32.000 0.000 32.000 0.000 40.000 16.568 40.000 40.000 16.568 40.000 -16.568 16.568 -40.000 ;
    LAYER M7 ;
    POLYGON -16.568 -40.000 -40.000 -16.568 -40.000 16.568 -16.568 40.000 0.000 40.000 0.000 32.000 -13.256 32.000 -32.000 13.256 -32.000 -13.256 -13.256 -32.000 13.256 -32.000 32.000 -13.256 32.000 13.256 13.256 32.000 0.000 32.000 0.000 40.000 16.568 40.000 40.000 16.568 40.000 -16.568 16.568 -40.000 ;
    LAYER M8 ;
    POLYGON -16.568 -40.000 -40.000 -16.568 -40.000 16.568 -16.568 40.000 0.000 40.000 0.000 32.000 -13.256 32.000 -32.000 13.256 -32.000 -13.256 -13.256 -32.000 13.256 -32.000 32.000 -13.256 32.000 13.256 13.256 32.000 0.000 32.000 0.000 40.000 16.568 40.000 40.000 16.568 40.000 -16.568 16.568 -40.000 ;
    LAYER M9 ;
    POLYGON -16.568 -40.000 -40.000 -16.568 -40.000 16.568 -16.568 40.000 0.000 40.000 0.000 32.000 -13.256 32.000 -32.000 13.256 -32.000 -13.256 -13.256 -32.000 13.256 -32.000 32.000 -13.256 32.000 13.256 13.256 32.000 0.000 32.000 0.000 40.000 16.568 40.000 40.000 16.568 40.000 -16.568 16.568 -40.000 ;
    LAYER M10 ;
    POLYGON -16.568 -40.000 -40.000 -16.568 -40.000 16.568 -16.568 40.000 0.000 40.000 0.000 32.000 -13.256 32.000 -32.000 13.256 -32.000 -13.256 -13.256 -32.000 13.256 -32.000 32.000 -13.256 32.000 13.256 13.256 32.000 0.000 32.000 0.000 40.000 16.568 40.000 40.000 16.568 40.000 -16.568 16.568 -40.000 ;
  END
END ALIGNMENT
