// //#############################################################################
// //# Function: Carry Save Adder (4:2) (aka 5:3)                                #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_csa42 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     input  b,
//     input  c,
//     input  d,
//     input  cin,
//     output sum,
//     output carry,
//     output cout
// );
// 
//     assign cout   = (a & b) | (b & c) | (a & c);
//     assign sumint = a ^ b ^ c;
//     assign sum    = cin ^ d ^ sumint;
//     assign carry  = (cin & d) | (cin & sumint) | (d & sumint);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_csa42.v:10.1-28.10" *)
module la_csa42 (
    a,
    b,
    c,
    d,
    cin,
    sum,
    carry,
    cout
);
  (* force_downto = 32'b00000000000000000000000000000001 *)
  (* src = "/home/pgadfort/.sc/cache/lambdapdk-v0.1.33/lambdapdk/gf180/libs/gf180mcu_fd_sc_mcu9t5v0/techmap/yosys/cells_adders.v:6.25-6.26" *)
  wire _00_;
  (* force_downto = 32'b00000000000000000000000000000001 *)
      (* src = "/home/pgadfort/.sc/cache/lambdapdk-v0.1.33/lambdapdk/gf180/libs/gf180mcu_fd_sc_mcu9t5v0/techmap/yosys/cells_adders.v:6.28-6.29" *)
  wire _01_;
  (* force_downto = 32'b00000000000000000000000000000001 *)
      (* src = "/home/pgadfort/.sc/cache/lambdapdk-v0.1.33/lambdapdk/gf180/libs/gf180mcu_fd_sc_mcu9t5v0/techmap/yosys/cells_adders.v:6.31-6.32" *)
  wire _02_;
  (* force_downto = 32'b00000000000000000000000000000001 *)
      (* src = "/home/pgadfort/.sc/cache/lambdapdk-v0.1.33/lambdapdk/gf180/libs/gf180mcu_fd_sc_mcu9t5v0/techmap/yosys/cells_adders.v:8.26-8.27" *)
  wire _03_;
  (* force_downto = 32'b00000000000000000000000000000001 *)
      (* src = "/home/pgadfort/.sc/cache/lambdapdk-v0.1.33/lambdapdk/gf180/libs/gf180mcu_fd_sc_mcu9t5v0/techmap/yosys/cells_adders.v:8.29-8.30" *)
  wire _04_;
  (* force_downto = 32'b00000000000000000000000000000001 *)
      (* src = "/home/pgadfort/.sc/cache/lambdapdk-v0.1.33/lambdapdk/gf180/libs/gf180mcu_fd_sc_mcu9t5v0/techmap/yosys/cells_adders.v:6.25-6.26" *)
  wire _05_;
  (* force_downto = 32'b00000000000000000000000000000001 *)
      (* src = "/home/pgadfort/.sc/cache/lambdapdk-v0.1.33/lambdapdk/gf180/libs/gf180mcu_fd_sc_mcu9t5v0/techmap/yosys/cells_adders.v:6.28-6.29" *)
  wire _06_;
  (* force_downto = 32'b00000000000000000000000000000001 *)
      (* src = "/home/pgadfort/.sc/cache/lambdapdk-v0.1.33/lambdapdk/gf180/libs/gf180mcu_fd_sc_mcu9t5v0/techmap/yosys/cells_adders.v:6.31-6.32" *)
  wire _07_;
  (* force_downto = 32'b00000000000000000000000000000001 *)
      (* src = "/home/pgadfort/.sc/cache/lambdapdk-v0.1.33/lambdapdk/gf180/libs/gf180mcu_fd_sc_mcu9t5v0/techmap/yosys/cells_adders.v:8.26-8.27" *)
  wire _08_;
  (* force_downto = 32'b00000000000000000000000000000001 *)
      (* src = "/home/pgadfort/.sc/cache/lambdapdk-v0.1.33/lambdapdk/gf180/libs/gf180mcu_fd_sc_mcu9t5v0/techmap/yosys/cells_adders.v:8.29-8.30" *)
  wire _09_;
  (* src = "inputs/la_csa42.v:13.12-13.13" *)
  input a;
  wire a;
  (* src = "inputs/la_csa42.v:14.12-14.13" *)
  input b;
  wire b;
  (* src = "inputs/la_csa42.v:15.12-15.13" *)
  input c;
  wire c;
  (* src = "inputs/la_csa42.v:19.12-19.17" *)
  output carry;
  wire carry;
  (* src = "inputs/la_csa42.v:17.12-17.15" *)
  input cin;
  wire cin;
  (* src = "inputs/la_csa42.v:20.12-20.16" *)
  output cout;
  wire cout;
  (* src = "inputs/la_csa42.v:16.12-16.13" *)
  input d;
  wire d;
  (* src = "inputs/la_csa42.v:18.12-18.15" *)
  output sum;
  wire sum;
  gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10_ (
      .I (a),
      .ZN(_00_)
  );
  gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11_ (
      .I (d),
      .ZN(_05_)
  );
  gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12_ (
      .I (b),
      .ZN(_01_)
  );
  gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13_ (
      .I (cin),
      .ZN(_06_)
  );
  gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14_ (
      .I (c),
      .ZN(_02_)
  );
  gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15_ (
      .I (_04_),
      .ZN(_07_)
  );
  gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16_ (
      .I (_09_),
      .ZN(sum)
  );
  gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17_ (
      .I (_03_),
      .ZN(cout)
  );
  gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18_ (
      .I (_08_),
      .ZN(carry)
  );
  (* module_not_derived = 32'b00000000000000000000000000000001 *)
      (* src = "/home/pgadfort/.sc/cache/lambdapdk-v0.1.33/lambdapdk/gf180/libs/gf180mcu_fd_sc_mcu9t5v0/techmap/yosys/cells_adders.v:42.41-44.12" *)
  gf180mcu_fd_sc_mcu9t5v0__addf_1 _19_ (
      .A (_00_),
      .B (_01_),
      .CI(_02_),
      .CO(_03_),
      .S (_04_)
  );
  (* module_not_derived = 32'b00000000000000000000000000000001 *)
      (* src = "/home/pgadfort/.sc/cache/lambdapdk-v0.1.33/lambdapdk/gf180/libs/gf180mcu_fd_sc_mcu9t5v0/techmap/yosys/cells_adders.v:42.41-44.12" *)
  gf180mcu_fd_sc_mcu9t5v0__addf_1 _20_ (
      .A (_05_),
      .B (_06_),
      .CI(_07_),
      .CO(_08_),
      .S (_09_)
  );
endmodule
