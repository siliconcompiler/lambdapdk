module \$_TBUF_ (input A, input E, output Y);
  gf180mcu_fd_sc_mcu7t5v0__bufz_1 _TECHMAP_REPLACE_ (
    .I(A),
    .Z(Y),
    .EN(E));
endmodule
