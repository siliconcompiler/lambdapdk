// //#############################################################################
// //# Function:  Positive edge-triggered static D-type flop-flop with async     #
// //#            active low preset.                                             #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_dffsq #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      clk,
//     input      nset,
//     output reg q
// );
// 
//     always @(posedge clk or negedge nset)
//         if (!nset) q <= 1'b1;
//         else q <= d;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_dffsq.v:11.1-24.10" *)
module la_dffsq (
    d,
    clk,
    nset,
    q
);
  (* src = "inputs/la_dffsq.v:15.16-15.19" *)
  input clk;
  wire clk;
  (* src = "inputs/la_dffsq.v:14.16-14.17" *)
  input d;
  wire d;
  (* src = "inputs/la_dffsq.v:16.16-16.20" *)
  input nset;
  wire nset;
  (* src = "inputs/la_dffsq.v:17.16-17.17" *)
  output q;
  wire q;
  (* src = "inputs/la_dffsq.v:20.5-22.21" *)
  sky130_fd_sc_hd__dfstp_2 _0_ (
      .CLK(clk),
      .D(d),
      .Q(q),
      .SET_B(nset)
  );
endmodule
