// //#############################################################################
// //# Function: Power isolation circuit                                         #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_isolo
//   #(parameter PROP = "DEFAULT")
//    (
//     input  iso, // isolation signal
//     input  in, // input
//     output out  // out = ~iso & in
//     );
// 
//    assign out = ~iso & in;
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_isolo(iso, in, out);
  wire _0_;
  input in;
  wire in;
  input iso;
  wire iso;
  output out;
  wire out;
  gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1_ (
    .I(iso),
    .ZN(_0_)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_2 _2_ (
    .A1(in),
    .A2(_0_),
    .Z(out)
  );
endmodule
