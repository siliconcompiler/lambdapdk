// //#############################################################################
// //# Function:  Positive edge-triggered static D-type flop-flop with async     #
// //#            active low preset and scan input.                              #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_sdffsq #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      si,
//     input      se,
//     input      clk,
//     input      nset,
//     output reg q
// );
// 
//   always @(posedge clk or negedge nset)
//     if (!nset) q <= 1'b1;
//     else q <= se ? si : d;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_sdffsq.v:11.1-26.10" *)
module la_sdffsq (
    d,
    si,
    se,
    clk,
    nset,
    q
);
  (* src = "inputs/la_sdffsq.v:22.3-24.27" *)
  wire _0_;
  (* unused_bits = "0" *)
  wire _1_;
  (* src = "inputs/la_sdffsq.v:17.16-17.19" *)
  input clk;
  wire clk;
  (* src = "inputs/la_sdffsq.v:14.16-14.17" *)
  input d;
  wire d;
  (* src = "inputs/la_sdffsq.v:18.16-18.20" *)
  input nset;
  wire nset;
  (* src = "inputs/la_sdffsq.v:19.16-19.17" *)
  output q;
  wire q;
  (* src = "inputs/la_sdffsq.v:16.16-16.18" *)
  input se;
  wire se;
  (* src = "inputs/la_sdffsq.v:15.16-15.18" *)
  input si;
  wire si;
  MUX2_X1 _2_ (
      .A(d),
      .B(si),
      .S(se),
      .Z(_0_)
  );
  (* src = "inputs/la_sdffsq.v:22.3-24.27" *)
  DFFS_X1 _3_ (
      .CK(clk),
      .D (_0_),
      .Q (q),
      .QN(_1_),
      .SN(nset)
  );
endmodule
