// //#############################################################################
// //# Function: Positive edge-triggered inverting static D-type flop-flop       #
// //#           with scan input.                                                #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_sdffqn #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      si,
//     input      se,
//     input      clk,
//     output reg qn
// );
// 
//     always @(posedge clk) qn <= se ? ~si : ~d;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
module la_sdffqn (
    d,
    si,
    se,
    clk,
    qn
);
  (* src = "generated" *)
  wire _0_;
  (* src = "generated" *)
  input clk;
  wire clk;
  (* src = "generated" *)
  input d;
  wire d;
  (* src = "generated" *)
  output qn;
  wire qn;
  (* src = "generated" *)
  input se;
  wire se;
  (* src = "generated" *)
  input si;
  wire si;
  sky130_fd_sc_hd__mux2i_2 _1_ (
      .A0(d),
      .A1(si),
      .S (se),
      .Y (_0_)
  );
  (* src = "generated" *)
  sky130_fd_sc_hd__dfxtp_1 _2_ (
      .CLK(clk),
      .D  (_0_),
      .Q  (qn)
  );
endmodule
