// //#############################################################################
// //# Function: Or-And (oa222) Gate                                             #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_oa222 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a0,
//     input  a1,
//     input  b0,
//     input  b1,
//     input  c0,
//     input  c1,
//     output z
// );
// 
//     assign z = (a0 | a1) & (b0 | b1) & (c0 | c1);
// 
// endmodule

/* Generated by Yosys 0.40+33 (git sha1 cd1fb8b15, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_oa222(a0, a1, b0, b1, c0, c1, z);
  wire _0_;
  wire _1_;
  wire _2_;
  input a0;
  wire a0;
  input a1;
  wire a1;
  input b0;
  wire b0;
  input b1;
  wire b1;
  input c0;
  wire c0;
  input c1;
  wire c1;
  output z;
  wire z;
  sg13g2_nor2_2 _3_ (
    .A(b1),
    .B(b0),
    .Y(_1_)
  );
  sg13g2_nor2_2 _4_ (
    .A(a1),
    .B(a0),
    .Y(_2_)
  );
  sg13g2_nor2_1 _5_ (
    .A(c1),
    .B(c0),
    .Y(_0_)
  );
  sg13g2_nor3_2 _6_ (
    .A(_1_),
    .B(_2_),
    .C(_0_),
    .Y(z)
  );
endmodule
