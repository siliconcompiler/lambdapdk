// //#############################################################################
// //# Function:  Positive edge-triggered static D-type flop-flop with async     #
// //#            active low preset.                                             #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_dffsq #(parameter PROP = "DEFAULT")   (
//     input      d,
//     input      clk,
//     input      nset,
//     output reg q
//     );
// 
//    always @ (posedge clk or negedge nset)
//      if(!nset)
//        q <= 1'b1;
//      else
//        q <= d;
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_dffsq(d, clk, nset, q);
  wire _0_;
  wire _1_;
  wire _2_;
  input clk;
  wire clk;
  input d;
  wire d;
  input nset;
  wire nset;
  output q;
  wire q;
  INVx2_ASAP7_75t_R _3_ (
    .A(nset),
    .Y(_1_)
  );
  INVx2_ASAP7_75t_R _4_ (
    .A(_0_),
    .Y(q)
  );
  ASYNC_DFFHx1_ASAP7_75t_R _5_ (
    .CLK(clk),
    .D(d),
    .QN(_0_),
    .RESET(_2_),
    .SET(_1_)
  );
  TIELOx1_ASAP7_75t_R _6_ (
    .L(_2_)
  );
endmodule
