// //#############################################################################
// //# Function: Carry Save Adder (4:2) (aka 5:3)                                #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_csa42 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     input  b,
//     input  c,
//     input  d,
//     input  cin,
//     output sum,
//     output carry,
//     output cout
// );
// 
//     assign cout   = (a & b) | (b & c) | (a & c);
//     assign sumint = a ^ b ^ c;
//     assign sum    = cin ^ d ^ sumint;
//     assign carry  = (cin & d) | (cin & sumint) | (d & sumint);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
module la_csa42 (
    a,
    b,
    c,
    d,
    cin,
    sum,
    carry,
    cout
);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  (* src = "generated" *)
  input a;
  wire a;
  (* src = "generated" *)
  input b;
  wire b;
  (* src = "generated" *)
  input c;
  wire c;
  (* src = "generated" *)
  output carry;
  wire carry;
  (* src = "generated" *)
  input cin;
  wire cin;
  (* src = "generated" *)
  output cout;
  wire cout;
  (* src = "generated" *)
  input d;
  wire d;
  (* src = "generated" *)
  output sum;
  wire sum;
  sg13g2_nor2_1 _08_ (
      .A(b),
      .B(a),
      .Y(_07_)
  );
  sg13g2_a21oi_2 _09_ (
      .A1(b),
      .A2(a),
      .B1(c),
      .Y (_00_)
  );
  sg13g2_nor2_2 _10_ (
      .A(_07_),
      .B(_00_),
      .Y(cout)
  );
  sg13g2_xor2_1 _11_ (
      .A(d),
      .B(cin),
      .X(_01_)
  );
  sg13g2_nand3_1 _12_ (
      .A(b),
      .B(a),
      .C(c),
      .Y(_02_)
  );
  sg13g2_nor3_1 _13_ (
      .A(b),
      .B(a),
      .C(c),
      .Y(_03_)
  );
  sg13g2_a21o_1 _14_ (
      .A1(cout),
      .A2(_02_),
      .B1(_03_),
      .X (_04_)
  );
  sg13g2_xnor2_1 _15_ (
      .A(_01_),
      .B(_04_),
      .Y(sum)
  );
  sg13g2_nand2_1 _16_ (
      .A(d),
      .B(cin),
      .Y(_05_)
  );
  sg13g2_nor2_1 _17_ (
      .A(d),
      .B(cin),
      .Y(_06_)
  );
  sg13g2_a21oi_1 _18_ (
      .A1(_05_),
      .A2(_04_),
      .B1(_06_),
      .Y (carry)
  );
endmodule
