// Source lambdapdk/sky130/libs/sky130io/lef/sky130_fd_io.lef

(* blackbox *)
module sky130_fd_io__overlay_vssd_lvc (
    inout AMUXBUS_A,
    inout AMUXBUS_B,
    inout VCCD,
    inout VCCHIB,
    inout VDDA,
    inout VDDIO,
    inout VDDIO_Q,
    inout VSSA,
    inout VSSD,
    inout VSSIO,
    inout VSSIO_Q,
    inout VSWITCH
);
endmodule

(* blackbox *)
module sky130_fd_io__overlay_vdda_hvc (
    inout AMUXBUS_A,
    inout AMUXBUS_B,
    inout VCCD,
    inout VCCHIB,
    inout VDDA,
    inout VDDIO,
    inout VDDIO_Q,
    inout VSSA,
    inout VSSD,
    inout VSSIO,
    inout VSSIO_Q,
    inout VSWITCH
);
endmodule

(* blackbox *)
module sky130_fd_io__overlay_vccd_hvc (
    inout AMUXBUS_A,
    inout AMUXBUS_B,
    inout VCCD,
    inout VCCHIB,
    inout VDDA,
    inout VDDIO,
    inout VDDIO_Q,
    inout VSSA,
    inout VSSD,
    inout VSSIO,
    inout VSSIO_Q,
    inout VSWITCH
);
endmodule

(* blackbox *)
module sky130_fd_io__corner_bus_overlay (
    inout AMUXBUS_A,
    inout AMUXBUS_B,
    inout VCCD,
    inout VCCHIB,
    inout VDDA,
    inout VDDIO,
    inout VDDIO_Q,
    inout VSSA,
    inout VSSD,
    inout VSSIO,
    inout VSSIO_Q,
    inout VSWITCH
);
endmodule

(* blackbox *)
module sky130_fd_io__top_ground_lvc_wpad (
    inout AMUXBUS_A,
    inout AMUXBUS_B,
    inout G_PAD,
    inout BDY2_B2B,
    inout DRN_LVC1,
    inout DRN_LVC2,
    inout G_CORE,
    inout OGC_LVC,
    inout SRC_BDY_LVC1,
    inout SRC_BDY_LVC2,
    inout VCCD,
    inout VCCHIB,
    inout VDDA,
    inout VDDIO,
    inout VDDIO_Q,
    inout VSSA,
    inout VSSD,
    inout VSSIO,
    inout VSSIO_Q,
    inout VSWITCH
);
endmodule

(* blackbox *)
module sky130_fd_io__overlay_vssa_hvc (
    inout AMUXBUS_A,
    inout AMUXBUS_B,
    inout VCCD,
    inout VCCHIB,
    inout VDDA,
    inout VDDIO,
    inout VDDIO_Q,
    inout VSSA,
    inout VSSD,
    inout VSSIO,
    inout VSSIO_Q,
    inout VSWITCH
);
endmodule

(* blackbox *)
module sky130_fd_io__top_power_hvc_wpadv2 (
    inout AMUXBUS_A,
    inout AMUXBUS_B,
    inout DRN_HVC,
    inout OGC_HVC,
    inout P_CORE,
    inout P_PAD,
    inout SRC_BDY_HVC,
    inout VCCD,
    inout VCCHIB,
    inout VDDA,
    inout VDDIO,
    inout VDDIO_Q,
    inout VSSA,
    inout VSSD,
    inout VSSIO,
    inout VSSIO_Q,
    inout VSWITCH
);
endmodule

(* blackbox *)
module sky130_fd_io__overlay_vccd_lvc (
    inout AMUXBUS_A,
    inout AMUXBUS_B,
    inout VCCD,
    inout VCCHIB,
    inout VDDA,
    inout VDDIO,
    inout VDDIO_Q,
    inout VSSA,
    inout VSSD,
    inout VSSIO,
    inout VSSIO_Q,
    inout VSWITCH
);
endmodule

(* blackbox *)
module sky130_fd_io__overlay_vssa_lvc (
    inout AMUXBUS_A,
    inout AMUXBUS_B,
    inout VCCD,
    inout VCCHIB,
    inout VDDA,
    inout VDDIO,
    inout VDDIO_Q,
    inout VSSA,
    inout VSSD,
    inout VSSIO,
    inout VSSIO_Q,
    inout VSWITCH
);
endmodule

(* blackbox *)
module sky130_fd_io__overlay_gpiov2 (
    inout AMUXBUS_A,
    inout AMUXBUS_B,
    inout PAD,
    inout VCCD,
    inout VCCHIB,
    inout VDDA,
    inout VDDIO,
    inout VDDIO_Q,
    inout VSSA,
    inout VSSD,
    inout VSSIO,
    inout VSSIO_Q,
    inout VSWITCH
);
endmodule

(* blackbox *)
module sky130_fd_io__overlay_vssio_lvc (
    inout AMUXBUS_A,
    inout AMUXBUS_B,
    inout VCCD,
    inout VCCHIB,
    inout VDDA,
    inout VDDIO,
    inout VDDIO_Q,
    inout VSSA,
    inout VSSD,
    inout VSSIO,
    inout VSSIO_Q,
    inout VSWITCH
);
endmodule

(* blackbox *)
module sky130_fd_io__overlay_vssio_hvc (
    inout AMUXBUS_A,
    inout AMUXBUS_B,
    inout VCCD,
    inout VCCHIB,
    inout VDDA,
    inout VDDIO,
    inout VDDIO_Q,
    inout VSSA,
    inout VSSD,
    inout VSSIO,
    inout VSSIO_Q,
    inout VSWITCH
);
endmodule

(* blackbox *)
module sky130_fd_io__overlay_vddio_lvc (
    inout AMUXBUS_A,
    inout AMUXBUS_B,
    inout VCCD,
    inout VCCHIB,
    inout VDDA,
    inout VDDIO,
    inout VDDIO_Q,
    inout VSSA,
    inout VSSD,
    inout VSSIO,
    inout VSSIO_Q,
    inout VSWITCH
);
endmodule

(* blackbox *)
module sky130_fd_io__top_power_lvc_wpad (
    inout AMUXBUS_A,
    inout AMUXBUS_B,
    inout P_PAD,
    inout BDY2_B2B,
    inout DRN_LVC1,
    inout DRN_LVC2,
    inout OGC_LVC,
    inout P_CORE,
    inout SRC_BDY_LVC1,
    inout SRC_BDY_LVC2,
    inout VCCD,
    inout VCCHIB,
    inout VDDA,
    inout VDDIO,
    inout VDDIO_Q,
    inout VSSA,
    inout VSSD,
    inout VSSIO,
    inout VSSIO_Q,
    inout VSWITCH
);
endmodule

(* blackbox *)
module sky130_fd_io__overlay_vddio_hvc (
    inout AMUXBUS_A,
    inout AMUXBUS_B,
    inout VCCD,
    inout VCCHIB,
    inout VDDA,
    inout VDDIO,
    inout VDDIO_Q,
    inout VSSA,
    inout VSSD,
    inout VSSIO,
    inout VSSIO_Q,
    inout VSWITCH
);
endmodule

(* blackbox *)
module sky130_fd_io__top_xres4v2 (
    inout AMUXBUS_A,
    inout AMUXBUS_B,
    input DISABLE_PULLUP_H,
    input ENABLE_H,
    input ENABLE_VDDIO,
    input EN_VDDIO_SIG_H,
    input FILT_IN_H,
    input INP_SEL_H,
    inout PAD,
    inout PAD_A_ESD_H,
    inout PULLUP_H,
    output TIE_HI_ESD,
    output TIE_LO_ESD,
    inout TIE_WEAK_HI_H,
    output XRES_H_N,
    input VCCD,
    input VCCHIB,
    input VDDA,
    input VDDIO,
    input VDDIO_Q,
    input VSSA,
    input VSSD,
    input VSSIO,
    input VSSIO_Q,
    input VSWITCH
);
endmodule

(* blackbox *)
module sky130_fd_io__top_gpio_ovtv2 (
    inout AMUXBUS_A,
    inout AMUXBUS_B,
    input ANALOG_EN,
    input ANALOG_POL,
    input ANALOG_SEL,
    input ENABLE_H,
    input ENABLE_INP_H,
    input ENABLE_VDDA_H,
    input ENABLE_VDDIO,
    input ENABLE_VSWITCH_H,
    input HLD_H_N,
    input HLD_OVR,
    input HYS_TRIM,
    output IN,
    input INP_DIS,
    output IN_H,
    input OE_N,
    input OUT,
    inout PAD,
    inout PAD_A_ESD_0_H,
    inout PAD_A_ESD_1_H,
    inout PAD_A_NOESD_H,
    input SLOW,
    output TIE_HI_ESD,
    output TIE_LO_ESD,
    input VINREF,
    input VTRIP_SEL,
    inout VCCD,
    inout VCCHIB,
    inout VDDA,
    inout VDDIO,
    inout VDDIO_Q,
    inout VSSA,
    inout VSSD,
    inout VSSIO,
    inout VSSIO_Q,
    inout VSWITCH,
    input [2:0] DM,
    input [1:0] IB_MODE_SEL,
    input [1:0] SLEW_CTL
);
endmodule

(* blackbox *)
module sky130_fd_io__overlay_vdda_lvc (
    inout AMUXBUS_A,
    inout AMUXBUS_B,
    inout VCCD,
    inout VCCHIB,
    inout VDDA,
    inout VDDIO,
    inout VDDIO_Q,
    inout VSSA,
    inout VSSD,
    inout VSSIO,
    inout VSSIO_Q,
    inout VSWITCH
);
endmodule

(* blackbox *)
module sky130_fd_io__overlay_vssd_hvc (
    inout AMUXBUS_A,
    inout AMUXBUS_B,
    inout VCCD,
    inout VCCHIB,
    inout VDDA,
    inout VDDIO,
    inout VDDIO_Q,
    inout VSSA,
    inout VSSD,
    inout VSSIO,
    inout VSSIO_Q,
    inout VSWITCH
);
endmodule

(* blackbox *)
module sky130_fd_io__top_gpiov2 (
    inout AMUXBUS_A,
    inout AMUXBUS_B,
    input ANALOG_EN,
    input ANALOG_POL,
    input ANALOG_SEL,
    input ENABLE_H,
    input ENABLE_INP_H,
    input ENABLE_VDDA_H,
    input ENABLE_VDDIO,
    input ENABLE_VSWITCH_H,
    input HLD_H_N,
    input HLD_OVR,
    input IB_MODE_SEL,
    output IN,
    input INP_DIS,
    output IN_H,
    input OE_N,
    input OUT,
    inout PAD,
    inout PAD_A_ESD_0_H,
    inout PAD_A_ESD_1_H,
    inout PAD_A_NOESD_H,
    input SLOW,
    output TIE_HI_ESD,
    output TIE_LO_ESD,
    input VTRIP_SEL,
    inout VCCD,
    inout VCCHIB,
    inout VDDA,
    inout VDDIO,
    inout VDDIO_Q,
    inout VSSA,
    inout VSSD,
    inout VSSIO,
    inout VSSIO_Q,
    inout VSWITCH,
    input [2:0] DM
);
endmodule

(* blackbox *)
module sky130_fd_io__top_ground_hvc_wpad (
    inout AMUXBUS_A,
    inout AMUXBUS_B,
    inout G_PAD,
    inout DRN_HVC,
    inout G_CORE,
    inout OGC_HVC,
    inout SRC_BDY_HVC,
    inout VCCD,
    inout VCCHIB,
    inout VDDA,
    inout VDDIO,
    inout VDDIO_Q,
    inout VSSA,
    inout VSSD,
    inout VSSIO,
    inout VSSIO_Q,
    inout VSWITCH
);
endmodule
