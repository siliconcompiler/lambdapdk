// //#############################################################################
// //# Function: Positive edge-triggered inverting static D-type flop-flop       #
// //#           with scan input.                                                #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_sdffqn #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      si,
//     input      se,
//     input      clk,
//     output reg qn
// );
// 
//     always @(posedge clk) qn <= se ? ~si : ~d;
// 
// endmodule

/* Generated by Yosys 0.40 (git sha1 a1bb0255d, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_sdffqn(d, si, se, clk, qn);
  wire _0_;
  wire _1_;
  wire _2_;
  wire _3_;
  input clk;
  wire clk;
  input d;
  wire d;
  output qn;
  wire qn;
  input se;
  wire se;
  input si;
  wire si;
  INVx1_ASAP7_75t_L _4_ (
    .A(si),
    .Y(_2_)
  );
  NOR2x1_ASAP7_75t_L _5_ (
    .A(d),
    .B(se),
    .Y(_3_)
  );
  AO21x1_ASAP7_75t_L _6_ (
    .A1(_2_),
    .A2(se),
    .B(_3_),
    .Y(_0_)
  );
  INVx1_ASAP7_75t_L _7_ (
    .A(_1_),
    .Y(qn)
  );
  DFFHQNx1_ASAP7_75t_L _8_ (
    .CLK(clk),
    .D(_0_),
    .QN(_1_)
  );
endmodule
