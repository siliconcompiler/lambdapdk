// //#############################################################################
// //# Function: Dual data rate input buffer                                     #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_iddr #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      clk,      // clock
//     input      in,       // data input sampled on both edges of clock
//     output reg outrise,  // rising edge sample
//     output reg outfall   // falling edge sample
// );
// 
//     // Negedge Sample
//     always @(negedge clk) outfall <= in;
// 
//     // Posedge Sample
//     reg inrise;
//     always @(posedge clk) inrise <= in;
// 
//     // Posedge Latch (for hold)
//     always @(clk or inrise) if (~clk) outrise <= inrise;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
(* keep_hierarchy *)
module la_iddr (
    clk,
    in,
    outrise,
    outfall
);
  wire _0_;
  (* src = "generated" *)
  input clk;
  wire clk;
  (* src = "generated" *)
  input in;
  wire in;
  (* src = "generated" *)
  wire inrise;
  (* src = "generated" *)
  output outfall;
  wire outfall;
  (* src = "generated" *)
  output outrise;
  wire outrise;
  sky130_fd_sc_hd__inv_2 _1_ (
      .A(clk),
      .Y(_0_)
  );
  (* module_not_derived = 32'b00000000000000000000000000000001 *) (* src = "generated" *)
  sky130_fd_sc_hd__dlxtn_1 _2_ (
      .D(inrise),
      .GATE_N(clk),
      .Q(outrise)
  );
  (* src = "generated" *)
  sky130_fd_sc_hd__dfxtp_1 _3_ (
      .CLK(clk),
      .D  (in),
      .Q  (inrise)
  );
  (* src = "generated" *)
  sky130_fd_sc_hd__dfxtp_1 _4_ (
      .CLK(_0_),
      .D  (in),
      .Q  (outfall)
  );
endmodule
