// //#############################################################################
// //# Function: Carry Save Adder (3:2)                                          #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_csa32 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     input  b,
//     input  c,
//     output sum,
//     output carry
// );
// 
//     assign sum   = a ^ b ^ c;
//     assign carry = (a & b) | (b & c) | (c & a);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_csa32.v:10.1-23.10" *)
module la_csa32 (
    a,
    b,
    c,
    sum,
    carry
);
  wire _0_;
  wire _1_;
  wire _2_;
  (* src = "inputs/la_csa32.v:13.12-13.13" *)
  input a;
  wire a;
  (* src = "inputs/la_csa32.v:14.12-14.13" *)
  input b;
  wire b;
  (* src = "inputs/la_csa32.v:15.12-15.13" *)
  input c;
  wire c;
  (* src = "inputs/la_csa32.v:17.12-17.17" *)
  output carry;
  wire carry;
  (* src = "inputs/la_csa32.v:16.12-16.15" *)
  output sum;
  wire sum;
  sky130_fd_sc_hdll__xnor2_2 _3_ (
      .A(b),
      .B(c),
      .Y(_0_)
  );
  sky130_fd_sc_hdll__xnor2_2 _4_ (
      .A(a),
      .B(_0_),
      .Y(sum)
  );
  sky130_fd_sc_hdll__nand2_1 _5_ (
      .A(b),
      .B(c),
      .Y(_1_)
  );
  sky130_fd_sc_hdll__o21ai_1 _6_ (
      .A1(b),
      .A2(c),
      .B1(a),
      .Y (_2_)
  );
  sky130_fd_sc_hdll__nand2_1 _7_ (
      .A(_1_),
      .B(_2_),
      .Y(carry)
  );
endmodule
