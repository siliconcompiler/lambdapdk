// //#############################################################################
// //# Function: Positive edge-triggered inverting static D-type flop-flop       #
// //#           with scan input.                                                #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_sdffqn #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      si,
//     input      se,
//     input      clk,
//     output reg qn
// );
// 
//     always @(posedge clk) qn <= se ? ~si : ~d;
// 
// endmodule

/* Generated by Yosys 0.40+33 (git sha1 cd1fb8b15, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_sdffqn(d, si, se, clk, qn);
  wire _0_;
  wire _1_;
  wire _2_;
  wire _3_;
  input clk;
  wire clk;
  input d;
  wire d;
  output qn;
  wire qn;
  input se;
  wire se;
  input si;
  wire si;
  sg13g2_nand2b_1 _4_ (
    .A_N(si),
    .B(se),
    .Y(_1_)
  );
  sg13g2_o21ai_1 _5_ (
    .A1(d),
    .A2(se),
    .B1(_1_),
    .Y(_0_)
  );
  sg13g2_dfrbp_1 _6_ (
    .CLK(clk),
    .D(_0_),
    .Q(qn),
    .Q_N(_2_),
    .RESET_B(_3_)
  );
  sg13g2_tiehi _7_ (
    .L_HI(_3_)
  );
endmodule
