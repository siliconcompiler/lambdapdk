// //#############################################################################
// //# Function: And-Or-Inverter (aoi211) Gate                                   #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_aoi211 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a0,
//     input  a1,
//     input  b0,
//     input  c0,
//     output z
// );
// 
//     assign z = ~((a0 & a1) | b0 | c0);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_aoi211.v:10.1-22.10" *)
module la_aoi211 (
    a0,
    a1,
    b0,
    c0,
    z
);
  (* src = "inputs/la_aoi211.v:13.12-13.14" *)
  input a0;
  wire a0;
  (* src = "inputs/la_aoi211.v:14.12-14.14" *)
  input a1;
  wire a1;
  (* src = "inputs/la_aoi211.v:15.12-15.14" *)
  input b0;
  wire b0;
  (* src = "inputs/la_aoi211.v:16.12-16.14" *)
  input c0;
  wire c0;
  (* src = "inputs/la_aoi211.v:17.12-17.13" *)
  output z;
  wire z;
  gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _0_ (
      .A1(a1),
      .A2(a0),
      .B (b0),
      .C (c0),
      .ZN(z)
  );
endmodule
