// //#############################################################################
// //# Function: Dual data rate input buffer                                     #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_iddr #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      clk,      // clock
//     input      in,       // data input sampled on both edges of clock
//     output reg outrise,  // rising edge sample
//     output reg outfall   // falling edge sample
// );
// 
//   // Negedge Sample
//   always @(negedge clk) outfall <= in;
// 
//   // Posedge Sample
//   reg inrise;
//   always @(posedge clk) inrise <= in;
// 
//   // Posedge Latch (for hold)
//   always @(clk or inrise) if (~clk) outrise <= inrise;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_iddr.v:10.1-29.10" *)
module la_iddr (
    clk,
    in,
    outrise,
    outfall
);
  (* src = "inputs/la_iddr.v:27.3-27.55|/home/pgadfort/lambdapdk/lambdapdk/gf180/libs/gf180mcu_fd_sc_mcu7t5v0/techmap/yosys/cells_latch.v:12.12-12.14" *)
  wire _0_;
  (* src = "inputs/la_iddr.v:13.16-13.19" *)
  input clk;
  wire clk;
  (* src = "inputs/la_iddr.v:14.16-14.18" *)
  input in;
  wire in;
  (* src = "inputs/la_iddr.v:23.7-23.13" *)
  wire inrise;
  (* src = "inputs/la_iddr.v:16.16-16.23" *)
  output outfall;
  wire outfall;
  (* src = "inputs/la_iddr.v:15.16-15.23" *)
  output outrise;
  wire outrise;
  gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1_ (
      .I (clk),
      .ZN(_0_)
  );
  (* module_not_derived = 32'b00000000000000000000000000000001 *)
      (* src = "inputs/la_iddr.v:27.3-27.55|/home/pgadfort/lambdapdk/lambdapdk/gf180/libs/gf180mcu_fd_sc_mcu7t5v0/techmap/yosys/cells_latch.v:10.37-14.10" *)
  gf180mcu_fd_sc_mcu7t5v0__latq_1 _2_ (
      .D(inrise),
      .E(_0_),
      .Q(outrise)
  );
  (* src = "inputs/la_iddr.v:24.3-24.38" *)
  gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3_ (
      .CLK(clk),
      .D  (in),
      .Q  (inrise)
  );
  (* src = "inputs/la_iddr.v:20.3-20.39" *)
  gf180mcu_fd_sc_mcu7t5v0__dffnq_2 _4_ (
      .CLKN(clk),
      .D(in),
      .Q(outfall)
  );
endmodule
