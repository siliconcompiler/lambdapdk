// //#############################################################################
// //# Function: Tie High Cell                                                   #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_tiehi #(
//     parameter PROP = "DEFAULT"
// ) (
//     output z
// );
// 
//     assign z = 1'b1;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
(* keep_hierarchy *)
module la_tiehi (
    z
);
  (* src = "generated" *)
  output z;
  wire z;
  TIEHIx1_ASAP7_75t_R _0_ (.H(z));
endmodule
