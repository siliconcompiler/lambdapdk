// //#############################################################################
// //# Function: 4-Input Mux                                                     #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_mux4 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  d0,
//     input  d1,
//     input  d2,
//     input  d3,
//     input  s0,
//     input  s1,
//     output z
// );
// 
//     assign z = (d0 & ~s1 & ~s0) | (d1 & ~s1 & s0) | (d2 & s1 & ~s0) | (d3 & s1 & s0);
// 
// endmodule

/* Generated by Yosys 0.40 (git sha1 a1bb0255d, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_mux4(d0, d1, d2, d3, s0, s1, z);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  input d0;
  wire d0;
  input d1;
  wire d1;
  input d2;
  wire d2;
  input d3;
  wire d3;
  input s0;
  wire s0;
  input s1;
  wire s1;
  output z;
  wire z;
  INVx1_ASAP7_75t_R _06_ (
    .A(s0),
    .Y(_04_)
  );
  INVx1_ASAP7_75t_R _07_ (
    .A(s1),
    .Y(_05_)
  );
  OR2x4_ASAP7_75t_R _08_ (
    .A(d0),
    .B(s1),
    .Y(_00_)
  );
  OA21x2_ASAP7_75t_R _09_ (
    .A1(_05_),
    .A2(d2),
    .B(_00_),
    .Y(_01_)
  );
  OR2x2_ASAP7_75t_R _10_ (
    .A(s1),
    .B(d1),
    .Y(_02_)
  );
  OA211x2_ASAP7_75t_R _11_ (
    .A1(_05_),
    .A2(d3),
    .B(_02_),
    .C(s0),
    .Y(_03_)
  );
  AO21x1_ASAP7_75t_R _12_ (
    .A1(_04_),
    .A2(_01_),
    .B(_03_),
    .Y(z)
  );
endmodule
