// //#############################################################################
// //# Function: 2-Input one-hot mux                                             #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_dmux2 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  sel1,
//     input  sel0,
//     input  in1,
//     input  in0,
//     output out
// );
// 
//     assign out = (sel0 & in0) | (sel1 & in1);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_dmux2.v:10.1-22.10" *)
module la_dmux2 (
    sel1,
    sel0,
    in1,
    in0,
    out
);
  wire _0_;
  (* src = "inputs/la_dmux2.v:16.12-16.15" *)
  input in0;
  wire in0;
  (* src = "inputs/la_dmux2.v:15.12-15.15" *)
  input in1;
  wire in1;
  (* src = "inputs/la_dmux2.v:17.12-17.15" *)
  output out;
  wire out;
  (* src = "inputs/la_dmux2.v:14.12-14.16" *)
  input sel0;
  wire sel0;
  (* src = "inputs/la_dmux2.v:13.12-13.16" *)
  input sel1;
  wire sel1;
  gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _1_ (
      .A1(in0),
      .A2(sel0),
      .B1(in1),
      .B2(sel1),
      .ZN(_0_)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_2 _2_ (
      .I (_0_),
      .ZN(out)
  );
endmodule
