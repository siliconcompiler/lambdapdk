// //#############################################################################
// //# Function:  D-type active-low transparent latch                            #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_latnq #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      clk,
//     output reg q
// );
// 
//     always @(clk or d) if (~clk) q <= d;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_latnq.v:10.1-20.10" *)
module la_latnq (
    d,
    clk,
    q
);
  (* src = "inputs/la_latnq.v:14.16-14.19" *)
  input clk;
  wire clk;
  (* src = "inputs/la_latnq.v:13.16-13.17" *)
  input d;
  wire d;
  (* src = "inputs/la_latnq.v:15.16-15.17" *)
  output q;
  wire q;
  (* module_not_derived = 32'b00000000000000000000000000000001 *)
      (* src = "inputs/la_latnq.v:18.5-18.41|/home/pgadfort/.sc/cache/lambdapdk-v0.1.33/lambdapdk/asap7/libs/asap7sc7p5t_lvt/techmap/yosys/cells_latch.v:10.23-14.10" *)
  DLLx1_ASAP7_75t_L _0_ (
      .CLK(clk),
      .D  (d),
      .Q  (q)
  );
endmodule
