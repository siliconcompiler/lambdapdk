// //#############################################################################
// //# Function: Power isolation circuit                                         #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_isohi #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  iso,  // isolation signal
//     input  in,   // input
//     output out   // out = iso | in
// );
// 
//   assign out = iso | in;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_isohi.v:10.1-20.10" *)
module la_isohi (
    iso,
    in,
    out
);
  (* src = "inputs/la_isohi.v:14.12-14.14" *)
  input in;
  wire in;
  (* src = "inputs/la_isohi.v:13.12-13.15" *)
  input iso;
  wire iso;
  (* src = "inputs/la_isohi.v:15.12-15.15" *)
  output out;
  wire out;
  OR2x2_ASAP7_75t_R _0_ (
      .A(in),
      .B(iso),
      .Y(out)
  );
endmodule
