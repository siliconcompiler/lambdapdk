/*****************************************************************************
 * Function: IO supply cell (vdda)
 * Copyright: Lambda Project Authors. All rights Reserved.
 * License:  MIT (see LICENSE file in Lambda repository)
 *
 * Docs:
 *
 *
 ****************************************************************************/
(* keep_hierarchy *)
module la_iovdda #(
    parameter PROP  = "DEFAULT",  // cell type
    parameter SIDE  = "NO",       // "NO", "SO", "EA", "WE"
    parameter RINGW = 8           // width of io ring
) (
    inout             vdd,    // core supply
    inout             vss,    // core ground
    inout             vddio,  // io supply
    inout             vssio,  // io ground
    inout [RINGW-1:0] ioring  // generic io-ring interface
);

  sg13g2_IOPadVdd iovdd (
    .iovdd(vddio),
    .iovss(vssio),
    .vdd(vdd),
    .vss(vss)
  );

endmodule
