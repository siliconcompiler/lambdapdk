// //#############################################################################
// //# Function: Positive edge-triggered inverting static D-type flop-flop       #
// //#           with scan input.                                                #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_sdffqn #(parameter PROP = "DEFAULT")   (
//     input      d,
//     input      si,
//     input      se,
//     input      clk,
//     output reg qn
//     );
// 
//    always @ (posedge clk)
//      qn <= se ? ~si : ~d;
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_sdffqn(d, si, se, clk, qn);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  input clk;
  wire clk;
  input d;
  wire d;
  output qn;
  wire qn;
  input se;
  wire se;
  input si;
  wire si;
  INVx2_ASAP7_75t_R _05_ (
    .A(si),
    .Y(_04_)
  );
  NOR2x1_ASAP7_75t_R _06_ (
    .A(d),
    .B(se),
    .Y(_03_)
  );
  AO21x1_ASAP7_75t_R _07_ (
    .A1(_04_),
    .A2(se),
    .B(_03_),
    .Y(_00_)
  );
  INVx2_ASAP7_75t_R _08_ (
    .A(clk),
    .Y(_02_)
  );
  INVx2_ASAP7_75t_R _09_ (
    .A(_01_),
    .Y(qn)
  );
  DFFLQNx2_ASAP7_75t_R _10_ (
    .CLK(_02_),
    .D(_00_),
    .QN(_01_)
  );
endmodule
