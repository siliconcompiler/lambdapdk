// //#############################################################################
// //# Function:  Positive edge-triggered static inverting D-type flop-flop with #
// //             async active low reset.                                        #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_dffrqn #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      clk,
//     input      nreset,
//     output reg qn
// );
// 
//     always @(posedge clk or negedge nreset)
//         if (!nreset) qn <= 1'b1;
//         else qn <= ~d;
// 
// endmodule

/* Generated by Yosys 0.40 (git sha1 a1bb0255d, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_dffrqn(d, clk, nreset, qn);
  wire _0_;
  wire _1_;
  wire _2_;
  input clk;
  wire clk;
  input d;
  wire d;
  input nreset;
  wire nreset;
  output qn;
  wire qn;
  INVx1_ASAP7_75t_L _3_ (
    .A(d),
    .Y(_0_)
  );
  INVx1_ASAP7_75t_L _4_ (
    .A(_1_),
    .Y(qn)
  );
  DFFASRHQNx1_ASAP7_75t_L _5_ (
    .CLK(clk),
    .D(_0_),
    .QN(_1_),
    .RESETN(nreset),
    .SETN(_2_)
  );
  TIEHIx1_ASAP7_75t_L _6_ (
    .H(_2_)
  );
endmodule
