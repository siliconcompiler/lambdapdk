// //#############################################################################
// //# Function:  D-type active-low transparent latch                            #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_latnq #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      clk,
//     output reg q
// );
// 
//     always @(clk or d) if (~clk) q <= d;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_latnq.v:10.1-20.10" *)
module la_latnq (
    d,
    clk,
    q
);
  (* src = "inputs/la_latnq.v:18.5-18.41|/home/pgadfort/.sc/cache/lambdapdk-v0.1.33/lambdapdk/ihp130/libs/sg13g2_stdcell/techmap/yosys/cells_latch.v:12.15-12.17" *)
  wire _0_;
  (* src = "inputs/la_latnq.v:14.16-14.19" *)
  input clk;
  wire clk;
  (* src = "inputs/la_latnq.v:13.16-13.17" *)
  input d;
  wire d;
  (* src = "inputs/la_latnq.v:15.16-15.17" *)
  output q;
  wire q;
  sg13g2_inv_2 _1_ (
      .A(clk),
      .Y(_0_)
  );
  (* module_not_derived = 32'b00000000000000000000000000000001 *)
      (* src = "inputs/la_latnq.v:18.5-18.41|/home/pgadfort/.sc/cache/lambdapdk-v0.1.33/lambdapdk/ihp130/libs/sg13g2_stdcell/techmap/yosys/cells_latch.v:10.19-14.10" *)
  sg13g2_dlhq_1 _2_ (
      .D(d),
      .GATE(_0_),
      .Q(q)
  );
endmodule
