// //#############################################################################
// //# Function: Tristate Buffer                                                 #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_tbuf #(parameter PROP = "DEFAULT")  (
//    input  a,
//    input  oe,
//    output z
//    );
// 
//    assign z = oe ? a : 1'bz;
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_tbuf(a, oe, z);
  input a;
  wire a;
  input oe;
  wire oe;
  output z;
  wire z;
  assign z = a;
endmodule
