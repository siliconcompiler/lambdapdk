// //#############################################################################
// //# Function: Positive edge-triggered inverting static D-type flop-flop       #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_dffqn #(parameter PROP = "DEFAULT")   (
//     input  	d,
//     input  	clk,
//     output reg  qn
//     );
// 
//    always @ (posedge clk)
//      qn <= ~d;
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_dffqn(d, clk, qn);
  wire _0_;
  wire _1_;
  wire _2_;
  input clk;
  wire clk;
  input d;
  wire d;
  output qn;
  wire qn;
  INVx2_ASAP7_75t_R _3_ (
    .A(d),
    .Y(_0_)
  );
  INVx2_ASAP7_75t_R _4_ (
    .A(clk),
    .Y(_2_)
  );
  INVx2_ASAP7_75t_R _5_ (
    .A(_1_),
    .Y(qn)
  );
  DFFLQNx2_ASAP7_75t_R _6_ (
    .CLK(_2_),
    .D(_0_),
    .QN(_1_)
  );
endmodule
