// //#############################################################################
// //# Function:  Positive edge-triggered static D-type flop-flop with async     #
// //#            active low preset.                                             #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_dffsq #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      clk,
//     input      nset,
//     output reg q
// );
// 
//     always @(posedge clk or negedge nset)
//         if (!nset) q <= 1'b1;
//         else q <= d;
// 
// endmodule

/* Generated by Yosys 0.40+33 (git sha1 cd1fb8b15, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_dffsq(d, clk, nset, q);
  wire _0_;
  wire _1_;
  input clk;
  wire clk;
  input d;
  wire d;
  input nset;
  wire nset;
  output q;
  wire q;
  sg13g2_inv_2 _2_ (
    .A(d),
    .Y(_0_)
  );
  sg13g2_dfrbp_1 _3_ (
    .CLK(clk),
    .D(_0_),
    .Q(_1_),
    .Q_N(q),
    .RESET_B(nset)
  );
endmodule
