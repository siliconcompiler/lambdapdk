// //#############################################################################
// //# Function:  Positive edge-triggered static inverting D-type flop-flop with #
// //             async active low set and scan input                            #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_sdffsqn #(parameter PROP = "DEFAULT")   (
//     input      d,
//     input      si,
//     input      se,
//     input      clk,
//     input      nset,
//     output reg qn
//     );
// 
//    always @ (posedge clk or negedge nset)
//      if(!nset)
//        qn <= 1'b0;
//      else
//        qn <= se ? ~si : ~d;
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_sdffsqn(d, si, se, clk, nset, qn);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  input clk;
  wire clk;
  input d;
  wire d;
  input nset;
  wire nset;
  output qn;
  wire qn;
  input se;
  wire se;
  input si;
  wire si;
  INVx2_ASAP7_75t_L _06_ (
    .A(si),
    .Y(_04_)
  );
  NOR2x1_ASAP7_75t_L _07_ (
    .A(d),
    .B(se),
    .Y(_03_)
  );
  AO21x1_ASAP7_75t_L _08_ (
    .A1(_04_),
    .A2(se),
    .B(_03_),
    .Y(_00_)
  );
  INVx2_ASAP7_75t_L _09_ (
    .A(nset),
    .Y(_02_)
  );
  INVx2_ASAP7_75t_L _10_ (
    .A(_01_),
    .Y(qn)
  );
  ASYNC_DFFHx1_ASAP7_75t_L _11_ (
    .CLK(clk),
    .D(_00_),
    .QN(_01_),
    .RESET(_02_),
    .SET(_05_)
  );
  TIELOx1_ASAP7_75t_L _12_ (
    .L(_05_)
  );
endmodule
