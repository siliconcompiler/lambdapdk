// //#############################################################################
// //# Function: Positive edge-triggered inverting static D-type flop-flop       #
// //#           with scan input.                                                #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_sdffqn #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      si,
//     input      se,
//     input      clk,
//     output reg qn
// );
// 
//     always @(posedge clk) qn <= se ? ~si : ~d;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
(* keep_hierarchy *)
module la_sdffqn (
    d,
    si,
    se,
    clk,
    qn
);
  (* src = "generated" *)
  wire _0_;
  wire _1_;
  (* unused_bits = "0" *)
  wire _2_;
  wire _3_;
  (* src = "generated" *)
  input clk;
  wire clk;
  (* src = "generated" *)
  input d;
  wire d;
  (* src = "generated" *)
  output qn;
  wire qn;
  (* src = "generated" *)
  input se;
  wire se;
  (* src = "generated" *)
  input si;
  wire si;
  sg13g2_nand2b_1 _4_ (
      .A_N(si),
      .B  (se),
      .Y  (_1_)
  );
  sg13g2_o21ai_1 _5_ (
      .A1(d),
      .A2(se),
      .B1(_1_),
      .Y (_0_)
  );
  (* src = "generated" *)
  sg13g2_dfrbp_1 _6_ (
      .CLK(clk),
      .D(_0_),
      .Q(qn),
      .Q_N(_2_),
      .RESET_B(_3_)
  );
  sg13g2_tiehi _7_ (.L_HI(_3_));
endmodule
