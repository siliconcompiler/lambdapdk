// //#############################################################################
// //# Function:  Positive edge-triggered static D-type flop-flop with async     #
// //#            active low reset and scan input                                #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_sdffrq #(parameter PROP = "DEFAULT")   (
//     input      d,
//     input      si,
//     input      se,
//     input      clk,
//     input      nreset,
//     output reg q
//     );
// 
//    always @ (posedge clk or negedge nreset)
//      if(!nreset)
//        q <= 1'b0;
//      else
//        q <= se ? si : d;
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_sdffrq(d, si, se, clk, nreset, q);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  input clk;
  wire clk;
  input d;
  wire d;
  input nreset;
  wire nreset;
  output q;
  wire q;
  input se;
  wire se;
  input si;
  wire si;
  INVx2_ASAP7_75t_SL _06_ (
    .A(se),
    .Y(_04_)
  );
  AND2x4_ASAP7_75t_SL _07_ (
    .A(si),
    .B(se),
    .Y(_03_)
  );
  AO21x1_ASAP7_75t_SL _08_ (
    .A1(d),
    .A2(_04_),
    .B(_03_),
    .Y(_00_)
  );
  INVx2_ASAP7_75t_SL _09_ (
    .A(nreset),
    .Y(_02_)
  );
  INVx2_ASAP7_75t_SL _10_ (
    .A(_01_),
    .Y(q)
  );
  ASYNC_DFFHx1_ASAP7_75t_SL _11_ (
    .CLK(clk),
    .D(_00_),
    .QN(_01_),
    .RESET(_02_),
    .SET(_05_)
  );
  TIELOx1_ASAP7_75t_SL _12_ (
    .L(_05_)
  );
endmodule
