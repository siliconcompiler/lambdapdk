// //#############################################################################
// //# Function:  Positive edge-triggered static D-type flop-flop with async     #
// //#            active low preset.                                             #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_dffsq #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      clk,
//     input      nset,
//     output reg q
// );
// 
//     always @(posedge clk or negedge nset)
//         if (!nset) q <= 1'b1;
//         else q <= d;
// 
// endmodule

/* Generated by Yosys 0.40 (git sha1 a1bb0255d, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_dffsq(d, clk, nset, q);
  wire _0_;
  wire _1_;
  input clk;
  wire clk;
  input d;
  wire d;
  input nset;
  wire nset;
  output q;
  wire q;
  INVx1_ASAP7_75t_SL _2_ (
    .A(_0_),
    .Y(q)
  );
  DFFASRHQNx1_ASAP7_75t_SL _3_ (
    .CLK(clk),
    .D(d),
    .QN(_0_),
    .RESETN(nset),
    .SETN(_1_)
  );
  TIEHIx1_ASAP7_75t_SL _4_ (
    .H(_1_)
  );
endmodule
