// //#############################################################################
// //# Function: 4-Input one-hot mux                                             #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_dmux4 #(
//     parameter PROP = "DEFAULT"  // cell property
// ) (
//     input  sel3,
//     input  sel2,
//     input  sel1,
//     input  sel0,
//     input  in3,
//     input  in2,
//     input  in1,
//     input  in0,
//     output out
// );
// 
//     assign out = (sel0 & in0) | (sel1 & in1) | (sel2 & in2) | (sel3 & in3);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_dmux4.v:10.1-26.10" *)
module la_dmux4 (
    sel3,
    sel2,
    sel1,
    sel0,
    in3,
    in2,
    in1,
    in0,
    out
);
  wire _0_;
  wire _1_;
  (* src = "inputs/la_dmux4.v:20.12-20.15" *)
  input in0;
  wire in0;
  (* src = "inputs/la_dmux4.v:19.12-19.15" *)
  input in1;
  wire in1;
  (* src = "inputs/la_dmux4.v:18.12-18.15" *)
  input in2;
  wire in2;
  (* src = "inputs/la_dmux4.v:17.12-17.15" *)
  input in3;
  wire in3;
  (* src = "inputs/la_dmux4.v:21.12-21.15" *)
  output out;
  wire out;
  (* src = "inputs/la_dmux4.v:16.12-16.16" *)
  input sel0;
  wire sel0;
  (* src = "inputs/la_dmux4.v:15.12-15.16" *)
  input sel1;
  wire sel1;
  (* src = "inputs/la_dmux4.v:14.12-14.16" *)
  input sel2;
  wire sel2;
  (* src = "inputs/la_dmux4.v:13.12-13.16" *)
  input sel3;
  wire sel3;
  AO22x1_ASAP7_75t_SL _2_ (
      .A1(in0),
      .A2(sel0),
      .B1(in2),
      .B2(sel2),
      .Y (_0_)
  );
  AO22x1_ASAP7_75t_SL _3_ (
      .A1(in1),
      .A2(sel1),
      .B1(in3),
      .B2(sel3),
      .Y (_1_)
  );
  OR2x2_ASAP7_75t_SL _4_ (
      .A(_0_),
      .B(_1_),
      .Y(out)
  );
endmodule
