// //#############################################################################
// //# Function: Synchronizer with async reset                                   #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// module la_drsync #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  clk,    // clock
//     input  in,     // input data
//     input  nreset, // async active low reset
//     output out     // synchronized data
// );
// 
//     localparam STAGES = 2;
// 
//     reg [STAGES-1:0] shiftreg;
// 
//     always @(posedge clk or negedge nreset)
//         if (!nreset) shiftreg[STAGES-1:0] <= 'b0;
//         else shiftreg[STAGES-1:0] <= {shiftreg[STAGES-2:0], in};
// 
//     assign out = shiftreg[STAGES-1];
// 
// endmodule

/* Generated by Yosys 0.41 (git sha1 c1ad37779, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_drsync(clk, in, nreset, out);
  wire _0_;
  wire _1_;
  input clk;
  wire clk;
  input in;
  wire in;
  input nreset;
  wire nreset;
  output out;
  wire out;
  wire \shiftreg[0] ;
  DFFR_X1 _2_ (
    .CK(clk),
    .D(in),
    .Q(\shiftreg[0] ),
    .QN(_1_),
    .RN(nreset)
  );
  DFFR_X1 _3_ (
    .CK(clk),
    .D(\shiftreg[0] ),
    .Q(out),
    .QN(_0_),
    .RN(nreset)
  );
endmodule
