// //#############################################################################
// //# Function: Inverter                                                        #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_inv #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     output z
// );
// 
//     assign z = ~a;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
(* keep_hierarchy *)
module la_inv (
    a,
    z
);
  (* src = "generated" *)
  input a;
  wire a;
  (* src = "generated" *)
  output z;
  wire z;
  sky130_fd_sc_hd__inv_2 _0_ (
      .A(a),
      .Y(z)
  );
endmodule
