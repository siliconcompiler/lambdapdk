// //#############################################################################
// //# Function: Carry Save Adder (4:2) (aka 5:3)                                #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_csa42 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     input  b,
//     input  c,
//     input  d,
//     input  cin,
//     output sum,
//     output carry,
//     output cout
// );
// 
//   assign cout   = (a & b) | (b & c) | (a & c);
//   assign sumint = a ^ b ^ c;
//   assign sum    = cin ^ d ^ sumint;
//   assign carry  = (cin & d) | (cin & sumint) | (d & sumint);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_csa42.v:10.1-28.10" *)
module la_csa42 (
    a,
    b,
    c,
    d,
    cin,
    sum,
    carry,
    cout
);
  (* force_downto = 32'b00000000000000000000000000000001 *)
  (* src = "/home/pgadfort/lambdapdk/lambdapdk/sky130/libs/sky130hd/techmap/yosys/cells_adders.v:6.25-6.26" *)
  wire _00_;
  (* force_downto = 32'b00000000000000000000000000000001 *)
      (* src = "/home/pgadfort/lambdapdk/lambdapdk/sky130/libs/sky130hd/techmap/yosys/cells_adders.v:6.28-6.29" *)
  wire _01_;
  (* force_downto = 32'b00000000000000000000000000000001 *)
      (* src = "/home/pgadfort/lambdapdk/lambdapdk/sky130/libs/sky130hd/techmap/yosys/cells_adders.v:6.31-6.32" *)
  wire _02_;
  (* force_downto = 32'b00000000000000000000000000000001 *)
      (* src = "/home/pgadfort/lambdapdk/lambdapdk/sky130/libs/sky130hd/techmap/yosys/cells_adders.v:8.26-8.27" *)
  wire _03_;
  (* force_downto = 32'b00000000000000000000000000000001 *)
      (* src = "/home/pgadfort/lambdapdk/lambdapdk/sky130/libs/sky130hd/techmap/yosys/cells_adders.v:8.29-8.30" *)
  wire _04_;
  (* force_downto = 32'b00000000000000000000000000000001 *)
      (* src = "/home/pgadfort/lambdapdk/lambdapdk/sky130/libs/sky130hd/techmap/yosys/cells_adders.v:6.25-6.26" *)
  wire _05_;
  (* force_downto = 32'b00000000000000000000000000000001 *)
      (* src = "/home/pgadfort/lambdapdk/lambdapdk/sky130/libs/sky130hd/techmap/yosys/cells_adders.v:6.28-6.29" *)
  wire _06_;
  (* force_downto = 32'b00000000000000000000000000000001 *)
      (* src = "/home/pgadfort/lambdapdk/lambdapdk/sky130/libs/sky130hd/techmap/yosys/cells_adders.v:6.31-6.32" *)
  wire _07_;
  (* force_downto = 32'b00000000000000000000000000000001 *)
      (* src = "/home/pgadfort/lambdapdk/lambdapdk/sky130/libs/sky130hd/techmap/yosys/cells_adders.v:8.26-8.27" *)
  wire _08_;
  (* force_downto = 32'b00000000000000000000000000000001 *)
      (* src = "/home/pgadfort/lambdapdk/lambdapdk/sky130/libs/sky130hd/techmap/yosys/cells_adders.v:8.29-8.30" *)
  wire _09_;
  (* src = "inputs/la_csa42.v:13.12-13.13" *)
  input a;
  wire a;
  (* src = "inputs/la_csa42.v:14.12-14.13" *)
  input b;
  wire b;
  (* src = "inputs/la_csa42.v:15.12-15.13" *)
  input c;
  wire c;
  (* src = "inputs/la_csa42.v:19.12-19.17" *)
  output carry;
  wire carry;
  (* src = "inputs/la_csa42.v:17.12-17.15" *)
  input cin;
  wire cin;
  (* src = "inputs/la_csa42.v:20.12-20.16" *)
  output cout;
  wire cout;
  (* src = "inputs/la_csa42.v:16.12-16.13" *)
  input d;
  wire d;
  (* src = "inputs/la_csa42.v:18.12-18.15" *)
  output sum;
  wire sum;
  sky130_fd_sc_hd__inv_2 _10_ (
      .A(a),
      .Y(_00_)
  );
  sky130_fd_sc_hd__inv_2 _11_ (
      .A(d),
      .Y(_05_)
  );
  sky130_fd_sc_hd__inv_2 _12_ (
      .A(b),
      .Y(_01_)
  );
  sky130_fd_sc_hd__inv_2 _13_ (
      .A(cin),
      .Y(_06_)
  );
  sky130_fd_sc_hd__inv_2 _14_ (
      .A(c),
      .Y(_02_)
  );
  sky130_fd_sc_hd__inv_2 _15_ (
      .A(_04_),
      .Y(_07_)
  );
  sky130_fd_sc_hd__inv_2 _16_ (
      .A(_09_),
      .Y(sum)
  );
  sky130_fd_sc_hd__inv_2 _17_ (
      .A(_03_),
      .Y(cout)
  );
  sky130_fd_sc_hd__inv_2 _18_ (
      .A(_08_),
      .Y(carry)
  );
  (* module_not_derived = 32'b00000000000000000000000000000001 *)
      (* src = "/home/pgadfort/lambdapdk/lambdapdk/sky130/libs/sky130hd/techmap/yosys/cells_adders.v:42.31-44.12" *)
  sky130_fd_sc_hd__fa_1 _19_ (
      .A(_00_),
      .B(_01_),
      .CIN(_02_),
      .COUT(_03_),
      .SUM(_04_)
  );
  (* module_not_derived = 32'b00000000000000000000000000000001 *)
      (* src = "/home/pgadfort/lambdapdk/lambdapdk/sky130/libs/sky130hd/techmap/yosys/cells_adders.v:42.31-44.12" *)
  sky130_fd_sc_hd__fa_1 _20_ (
      .A(_05_),
      .B(_06_),
      .CIN(_07_),
      .COUT(_08_),
      .SUM(_09_)
  );
endmodule
