// //#############################################################################
// //# Function: Dual data rate input buffer                                     #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_iddr #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      clk,      // clock
//     input      in,       // data input sampled on both edges of clock
//     output reg outrise,  // rising edge sample
//     output reg outfall   // falling edge sample
// );
// 
//     // Negedge Sample
//     always @(negedge clk) outfall <= in;
// 
//     // Posedge Sample
//     reg inrise;
//     always @(posedge clk) inrise <= in;
// 
//     // Posedge Latch (for hold)
//     always @(clk or inrise) if (~clk) outrise <= inrise;
// 
// endmodule

/* Generated by Yosys 0.40 (git sha1 a1bb0255d, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_iddr(clk, in, outrise, outfall);
  wire _0_;
  wire _1_;
  input clk;
  wire clk;
  input in;
  wire in;
  wire inrise;
  output outfall;
  wire outfall;
  output outrise;
  wire outrise;
  INVx1_ASAP7_75t_SL _2_ (
    .A(_0_),
    .Y(outfall)
  );
  INVx1_ASAP7_75t_SL _3_ (
    .A(_1_),
    .Y(inrise)
  );
  DLLx1_ASAP7_75t_SL _4_ (
    .CLK(clk),
    .D(inrise),
    .Q(outrise)
  );
  DFFHQNx1_ASAP7_75t_SL _5_ (
    .CLK(clk),
    .D(in),
    .QN(_1_)
  );
  DFFLQNx1_ASAP7_75t_SL _6_ (
    .CLK(clk),
    .D(in),
    .QN(_0_)
  );
endmodule
