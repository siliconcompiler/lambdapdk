// //#############################################################################
// //# Function: Or-And-Inverter (oai221) Gate                                   #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_oai221 #(parameter PROP = "DEFAULT")   (
//     input  a0,
//     input  a1,
//     input  b0,
//     input  b1,
//     input  c0,
//     output z
//     );
// 
//    assign z = ~((a0 | a1) & (b0 | b1) & (c0));
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_oai221(a0, a1, b0, b1, c0, z);
  wire _0_;
  wire _1_;
  input a0;
  wire a0;
  input a1;
  wire a1;
  input b0;
  wire b0;
  input b1;
  wire b1;
  input c0;
  wire c0;
  output z;
  wire z;
  OR2x2_ASAP7_75t_SL _2_ (
    .A(a1),
    .B(a0),
    .Y(_0_)
  );
  OA21x2_ASAP7_75t_SL _3_ (
    .A1(b1),
    .A2(b0),
    .B(c0),
    .Y(_1_)
  );
  NAND2x1_ASAP7_75t_SL _4_ (
    .A(_0_),
    .B(_1_),
    .Y(z)
  );
endmodule
