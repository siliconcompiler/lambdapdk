// //#############################################################################
// //# Function:  Reset synchronizer (async assert, sync deassert)               #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_rsync
//   #(parameter PROP = "DEFAULT")
//    (
//     input  clk, // clock
//     input  nrst_in, // async reset input
//     output nrst_out // async assert, sync deassert reset
//    );
// 
//    localparam STAGES=2;
//    localparam RND = 1;
// 
//    reg [STAGES:0] sync_pipe;
//    integer        sync_delay;
// 
// `ifndef SYNTHESIS
//    always @ (posedge clk)
//      sync_delay <= {$random} % 2;
// `endif
// 
//    always @ (posedge clk or negedge nrst_in)
//      if(!nrst_in)
//        sync_pipe[STAGES:0] <= 'b0;
//      else
//        sync_pipe[STAGES:0] <= {sync_pipe[STAGES-1:0],1'b1};
// 
// `ifdef SYNTHESIS
//    assign nrst_out = sync_pipe[STAGES-1];
// `else
//    assign nrst_out = (|sync_delay & (|RND)) ? sync_pipe[STAGES] : sync_pipe[STAGES-1];
// `endif
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_rsync(clk, nrst_in, nrst_out);
  wire _0_;
  input clk;
  wire clk;
  input nrst_in;
  wire nrst_in;
  output nrst_out;
  wire nrst_out;
  wire \sync_pipe[0] ;
  gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _1_ (
    .CLK(clk),
    .D(_0_),
    .Q(\sync_pipe[0] ),
    .RN(nrst_in)
  );
  gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _2_ (
    .CLK(clk),
    .D(\sync_pipe[0] ),
    .Q(nrst_out),
    .RN(nrst_in)
  );
  gf180mcu_fd_sc_mcu7t5v0__tieh _3_ (
    .Z(_0_)
  );
endmodule
