// //#############################################################################
// //# Function: Non-inverting buffer with supplies                              #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_pwrbuf #(
//     parameter TARGET = "DEFAULT",  // "SIM"
//     parameter PROP   = "DEFAULT"
// ) (
//     input  vdd,
//     input  vss,
//     input  a,
//     output z
// );
// 
//     generate
//         if (TARGET == "SIM") assign z = ((vdd === 1'b1) && (vss === 1'b0)) ? a : 1'bX;
//         else assign z = a;
//     endgenerate
// 
// endmodule

/* Generated by Yosys 0.38+92 (git sha1 84116c9a3, x86_64-conda-linux-gnu-cc 11.2.0 -fvisibility-inlines-hidden -fmessage-length=0 -march=nocona -mtune=haswell -ftree-vectorize -fPIC -fstack-protector-strong -fno-plt -O2 -ffunction-sections -fdebug-prefix-map=/root/conda-eda/conda-eda/workdir/conda-env/conda-bld/yosys_1708682838165/work=/usr/local/src/conda/yosys-0.38_93_g84116c9a3 -fdebug-prefix-map=/user/projekt_pia/miniconda3/envs/sc=/usr/local/src/conda-prefix -fPIC -Os -fno-merge-constants) */

module la_pwrbuf(vdd, vss, a, z);
  input a;
  wire a;
  input vdd;
  wire vdd;
  input vss;
  wire vss;
  output z;
  wire z;
  assign z = a;
endmodule
