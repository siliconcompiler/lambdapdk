// //#############################################################################
// //# Function: 5-Input one-hot mux                                             #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_dmux5 #(
//     parameter PROP = "DEFAULT"  // cell property
// ) (
//     input  sel4,
//     input  sel3,
//     input  sel2,
//     input  sel1,
//     input  sel0,
//     input  in4,
//     input  in3,
//     input  in2,
//     input  in1,
//     input  in0,
//     output out
// );
// 
//     assign out = (sel0 & in0) | (sel1 & in1) | (sel2 & in2) | (sel3 & in3) | (sel4 & in4);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
(* keep_hierarchy *)
module la_dmux5 (
    sel4,
    sel3,
    sel2,
    sel1,
    sel0,
    in4,
    in3,
    in2,
    in1,
    in0,
    out
);
  wire _0_;
  wire _1_;
  (* src = "generated" *)
  input in0;
  wire in0;
  (* src = "generated" *)
  input in1;
  wire in1;
  (* src = "generated" *)
  input in2;
  wire in2;
  (* src = "generated" *)
  input in3;
  wire in3;
  (* src = "generated" *)
  input in4;
  wire in4;
  (* src = "generated" *)
  output out;
  wire out;
  (* src = "generated" *)
  input sel0;
  wire sel0;
  (* src = "generated" *)
  input sel1;
  wire sel1;
  (* src = "generated" *)
  input sel2;
  wire sel2;
  (* src = "generated" *)
  input sel3;
  wire sel3;
  (* src = "generated" *)
  input sel4;
  wire sel4;
  sky130_fd_sc_hdll__a22oi_1 _2_ (
      .A1(in0),
      .A2(sel0),
      .B1(in4),
      .B2(sel4),
      .Y (_0_)
  );
  sky130_fd_sc_hdll__a222oi_1 _3_ (
      .A1(in1),
      .A2(sel1),
      .B1(in2),
      .B2(sel2),
      .C1(in3),
      .C2(sel3),
      .Y (_1_)
  );
  sky130_fd_sc_hdll__nand2_1 _4_ (
      .A(_0_),
      .B(_1_),
      .Y(out)
  );
endmodule
