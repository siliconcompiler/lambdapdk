// //#############################################################################
// //# Function: 4 Input Nor Gate                                                #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_nor4 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     input  b,
//     input  c,
//     input  d,
//     output z
// );
// 
//     assign z = ~(a | b | c | d);
// 
// endmodule

/* Generated by Yosys 0.40 (git sha1 a1bb0255d, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_nor4(a, b, c, d, z);
  wire _0_;
  input a;
  wire a;
  input b;
  wire b;
  input c;
  wire c;
  input d;
  wire d;
  output z;
  wire z;
  OR4x1_ASAP7_75t_R _1_ (
    .A(b),
    .B(a),
    .C(c),
    .D(d),
    .Y(_0_)
  );
  INVx1_ASAP7_75t_R _2_ (
    .A(_0_),
    .Y(z)
  );
endmodule
