// //#############################################################################
// //# Function: And-Or (ao33) Gate                                              #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_ao33 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a0,
//     input  a1,
//     input  a2,
//     input  b0,
//     input  b1,
//     input  b2,
//     output z
// );
// 
//     assign z = (a0 & a1 & a2) | (b0 & b1 & b2);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_ao33.v:10.1-24.10" *)
module la_ao33 (
    a0,
    a1,
    a2,
    b0,
    b1,
    b2,
    z
);
  wire _0_;
  wire _1_;
  (* src = "inputs/la_ao33.v:13.12-13.14" *)
  input a0;
  wire a0;
  (* src = "inputs/la_ao33.v:14.12-14.14" *)
  input a1;
  wire a1;
  (* src = "inputs/la_ao33.v:15.12-15.14" *)
  input a2;
  wire a2;
  (* src = "inputs/la_ao33.v:16.12-16.14" *)
  input b0;
  wire b0;
  (* src = "inputs/la_ao33.v:17.12-17.14" *)
  input b1;
  wire b1;
  (* src = "inputs/la_ao33.v:18.12-18.14" *)
  input b2;
  wire b2;
  (* src = "inputs/la_ao33.v:19.12-19.13" *)
  output z;
  wire z;
  sky130_fd_sc_hdll__nand3_2 _2_ (
      .A(b2),
      .B(b1),
      .C(b0),
      .Y(_0_)
  );
  sky130_fd_sc_hdll__nand3_2 _3_ (
      .A(a1),
      .B(a0),
      .C(a2),
      .Y(_1_)
  );
  sky130_fd_sc_hdll__nand2_2 _4_ (
      .A(_0_),
      .B(_1_),
      .Y(z)
  );
endmodule
