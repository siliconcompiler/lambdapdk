// //#############################################################################
// //# Function: Synchronizer with async reset                                   #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// module la_drsync #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  clk,    // clock
//     input  in,     // input data
//     input  nreset, // async active low reset
//     output out     // synchronized data
// );
// 
//   localparam STAGES = 2;
// 
//   reg [STAGES-1:0] shiftreg;
// 
//   always @(posedge clk or negedge nreset)
//     if (!nreset) shiftreg[STAGES-1:0] <= 'b0;
//     else shiftreg[STAGES-1:0] <= {shiftreg[STAGES-2:0], in};
// 
//   assign out = shiftreg[STAGES-1];
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* dynports =  1  *)
(* top =  1  *)
(* src = "inputs/la_drsync.v:9.1-28.10" *)
module la_drsync (
    clk,
    in,
    nreset,
    out
);
  (* src = "inputs/la_drsync.v:12.12-12.15" *)
  input clk;
  wire clk;
  (* src = "inputs/la_drsync.v:13.12-13.14" *)
  input in;
  wire in;
  (* src = "inputs/la_drsync.v:14.12-14.18" *)
  input nreset;
  wire nreset;
  (* src = "inputs/la_drsync.v:15.12-15.15" *)
  output out;
  wire out;
  (* src = "inputs/la_drsync.v:20.20-20.28" *)
  wire \shiftreg[0] ;
  (* src = "inputs/la_drsync.v:22.3-24.61" *)
  sky130_fd_sc_hdll__dfrtp_1 _0_ (
      .CLK(clk),
      .D(in),
      .Q(\shiftreg[0] ),
      .RESET_B(nreset)
  );
  (* src = "inputs/la_drsync.v:22.3-24.61" *)
  sky130_fd_sc_hdll__dfrtp_1 _1_ (
      .CLK(clk),
      .D(\shiftreg[0] ),
      .Q(out),
      .RESET_B(nreset)
  );
endmodule
