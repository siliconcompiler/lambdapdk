// //#############################################################################
// //# Function:  Positive edge-triggered static inverting D-type flop-flop with #
// //             async active low set.                                          #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_dffsqn #(parameter PROP = "DEFAULT")   (
//     input d,
//     input clk,
//     input nset,
//     output reg  qn
//     );
// 
//    always @ (posedge clk or negedge nset)
//      if(!nset)
//        qn <= 1'b0;
//      else
//        qn <= ~d;
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_dffsqn(d, clk, nset, qn);
  wire _0_;
  wire _1_;
  wire _2_;
  wire _3_;
  input clk;
  wire clk;
  input d;
  wire d;
  input nset;
  wire nset;
  output qn;
  wire qn;
  INVx2_ASAP7_75t_SL _4_ (
    .A(d),
    .Y(_0_)
  );
  INVx2_ASAP7_75t_SL _5_ (
    .A(nset),
    .Y(_2_)
  );
  INVx2_ASAP7_75t_SL _6_ (
    .A(_1_),
    .Y(qn)
  );
  ASYNC_DFFHx1_ASAP7_75t_SL _7_ (
    .CLK(clk),
    .D(_0_),
    .QN(_1_),
    .RESET(_2_),
    .SET(_3_)
  );
  TIELOx1_ASAP7_75t_SL _8_ (
    .L(_3_)
  );
endmodule
