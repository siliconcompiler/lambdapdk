// //#############################################################################
// //# Function: Positive edge-triggered static D-type flop-flop with scan input #
// //#                                                                           #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_sdffq #(parameter PROP = "DEFAULT")   (
//     input      d,
//     input      si,
//     input      se,
//     input      clk,
//     output reg q
//     );
// 
//    always @ (posedge clk)
//        q <= se ? si : d;
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_sdffq(d, si, se, clk, q);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  input clk;
  wire clk;
  input d;
  wire d;
  output q;
  wire q;
  input se;
  wire se;
  input si;
  wire si;
  INVx2_ASAP7_75t_SL _05_ (
    .A(se),
    .Y(_04_)
  );
  AND2x4_ASAP7_75t_SL _06_ (
    .A(si),
    .B(se),
    .Y(_03_)
  );
  AO21x1_ASAP7_75t_SL _07_ (
    .A1(d),
    .A2(_04_),
    .B(_03_),
    .Y(_00_)
  );
  INVx2_ASAP7_75t_SL _08_ (
    .A(clk),
    .Y(_02_)
  );
  INVx2_ASAP7_75t_SL _09_ (
    .A(_01_),
    .Y(q)
  );
  DFFLQNx2_ASAP7_75t_SL _10_ (
    .CLK(_02_),
    .D(_00_),
    .QN(_01_)
  );
endmodule
