// //#############################################################################
// //# Function: Carry Save Adder (3:2)                                          #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_csa32 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     input  b,
//     input  c,
//     output sum,
//     output carry
// );
// 
//     assign sum   = a ^ b ^ c;
//     assign carry = (a & b) | (b & c) | (c & a);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_csa32.v:10.1-23.10" *)
module la_csa32 (
    a,
    b,
    c,
    sum,
    carry
);
  (* src = "/home/pgadfort/.sc/cache/lambdapdk-v0.1.33/lambdapdk/asap7/libs/asap7sc7p5t_slvt/techmap/yosys/cells_adders.v:10.22-10.24" *)
  wire _0_;
  (* src = "/home/pgadfort/.sc/cache/lambdapdk-v0.1.33/lambdapdk/asap7/libs/asap7sc7p5t_slvt/techmap/yosys/cells_adders.v:10.26-10.28" *)
  wire _1_;
  (* src = "inputs/la_csa32.v:13.12-13.13" *)
  input a;
  wire a;
  (* src = "inputs/la_csa32.v:14.12-14.13" *)
  input b;
  wire b;
  (* src = "inputs/la_csa32.v:15.12-15.13" *)
  input c;
  wire c;
  (* src = "inputs/la_csa32.v:17.12-17.17" *)
  output carry;
  wire carry;
  (* src = "inputs/la_csa32.v:16.12-16.15" *)
  output sum;
  wire sum;
  INVx2_ASAP7_75t_SL _2_ (
      .A(_0_),
      .Y(carry)
  );
  INVx2_ASAP7_75t_SL _3_ (
      .A(_1_),
      .Y(sum)
  );
  (* module_not_derived = 32'b00000000000000000000000000000001 *)
      (* src = "/home/pgadfort/.sc/cache/lambdapdk-v0.1.33/lambdapdk/asap7/libs/asap7sc7p5t_slvt/techmap/yosys/cells_adders.v:44.27-46.12" *)
  FAx1_ASAP7_75t_SL _4_ (
      .A  (a),
      .B  (b),
      .CI (c),
      .CON(_0_),
      .SN (_1_)
  );
endmodule
