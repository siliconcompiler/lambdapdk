// //#############################################################################
// //# Function:  Positive edge-triggered static inverting D-type flop-flop with #
// //             async active low reset.                                        #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_dffrqn #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      clk,
//     input      nreset,
//     output reg qn
// );
// 
//     always @(posedge clk or negedge nreset)
//         if (!nreset) qn <= 1'b1;
//         else qn <= ~d;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_dffrqn.v:11.1-24.10" *)
module la_dffrqn (
    d,
    clk,
    nreset,
    qn
);
  (* src = "inputs/la_dffrqn.v:20.5-22.23" *)
  wire _0_;
  (* src = "inputs/la_dffrqn.v:15.16-15.19" *)
  input clk;
  wire clk;
  (* src = "inputs/la_dffrqn.v:14.16-14.17" *)
  input d;
  wire d;
  (* src = "inputs/la_dffrqn.v:16.16-16.22" *)
  input nreset;
  wire nreset;
  (* src = "inputs/la_dffrqn.v:17.16-17.18" *)
  output qn;
  wire qn;
  gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1_ (
      .I (d),
      .ZN(_0_)
  );
  (* src = "inputs/la_dffrqn.v:20.5-22.23" *)
  gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 _2_ (
      .CLK(clk),
      .D(_0_),
      .Q(qn),
      .SETN(nreset)
  );
endmodule
