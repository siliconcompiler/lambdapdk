
//Solution to the short was found at the end of a conversation thread at this
//link:
//https://groups.google.com/g/comp.lang.verilog/c/b3-6XMA8KA4

module la_pt (
    .io1(a),
    .io2(a)
);
    inout wire a;
endmodule  // la_pt
