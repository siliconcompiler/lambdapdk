// //#############################################################################
// //# Function: 3-Input one-hot mux                                             #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_dmux3 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  sel0,
//     input  sel1,
//     input  sel2,
//     input  in0,
//     input  in1,
//     input  in2,
//     output out
// );
// 
//     assign out = (sel0 & in0) | (sel1 & in1) | (sel2 & in2);
// 
// endmodule

/* Generated by Yosys 0.38+92 (git sha1 84116c9a3, x86_64-conda-linux-gnu-cc 11.2.0 -fvisibility-inlines-hidden -fmessage-length=0 -march=nocona -mtune=haswell -ftree-vectorize -fPIC -fstack-protector-strong -fno-plt -O2 -ffunction-sections -fdebug-prefix-map=/root/conda-eda/conda-eda/workdir/conda-env/conda-bld/yosys_1708682838165/work=/usr/local/src/conda/yosys-0.38_93_g84116c9a3 -fdebug-prefix-map=/user/projekt_pia/miniconda3/envs/sc=/usr/local/src/conda-prefix -fPIC -Os -fno-merge-constants) */

module la_dmux3(sel0, sel1, sel2, in0, in1, in2, out);
  wire _0_;
  input in0;
  wire in0;
  input in1;
  wire in1;
  input in2;
  wire in2;
  output out;
  wire out;
  input sel0;
  wire sel0;
  input sel1;
  wire sel1;
  input sel2;
  wire sel2;
  sky130_fd_sc_hdll__a222oi_1 _1_ (
    .A1(in0),
    .A2(sel0),
    .B1(in1),
    .B2(sel1),
    .C1(in2),
    .C2(sel2),
    .Y(_0_)
  );
  sky130_fd_sc_hdll__inv_1 _2_ (
    .A(_0_),
    .Y(out)
  );
endmodule
