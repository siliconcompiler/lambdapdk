# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

#=====================================
# Revision: 1.1
#=====================================

VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS   1000 ;
END UNITS

MANUFACTURINGGRID   0.005 ;



MACRO gf180mcu_fd_ip_sram__sram512x8m8wm1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_fd_ip_sram__sram512x8m8wm1 0 0 ;
  SIZE 431.86 BY 484.88 ;
  SYMMETRY X Y R90 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.9976 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 171.215 0 172.335 1 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.9976 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 162.76 0 163.88 1 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.9976 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 154.295 0 155.415 1 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.9976 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 281.325 0 282.445 1 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.9976 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 275.82 0 276.94 1 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.9976 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 272.085 0 273.205 1 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.9976 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 268.86 0 269.98 1 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.9976 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 148.525 0 149.645 1 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.9976 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 145.03 0 146.15 1 ;
    END
  END A[8]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.9976 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 251.71 0 252.83 1 ;
    END
  END CEN
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
      ANTENNAGATEAREA 44.7066 LAYER Metal3 ;
      ANTENNAGATEAREA 2.868 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 139.68 0 140.8 1 ;
    END
  END CLK
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
      ANTENNAGATEAREA 1.152 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 9.32 0 10.44 1 ;
    END
  END D[0]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
      ANTENNAGATEAREA 1.152 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 61.03 0 62.15 1 ;
    END
  END D[1]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
      ANTENNAGATEAREA 1.152 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 67.27 0 68.39 1 ;
    END
  END D[2]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
      ANTENNAGATEAREA 1.152 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 118.975 0 120.095 1 ;
    END
  END D[3]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
      ANTENNAGATEAREA 1.152 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 307.235 0 308.355 1 ;
    END
  END D[4]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
      ANTENNAGATEAREA 1.152 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 358.91 0 360.03 1 ;
    END
  END D[5]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
      ANTENNAGATEAREA 1.152 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 365.15 0 366.27 1 ;
    END
  END D[6]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
      ANTENNAGATEAREA 1.152 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 416.86 0 417.98 1 ;
    END
  END D[7]
  PIN GWEN
    DIRECTION INPUT ;
    USE SIGNAL ;
      ANTENNAGATEAREA 14.466 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 202.94 0 204.06 1 ;
    END
  END GWEN
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.328 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 16.9 0 18.02 1 ;
    END
  END Q[0]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.328 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 57.665 0 58.785 1 ;
    END
  END Q[1]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.328 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 70.635 0 71.755 1 ;
    END
  END Q[2]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.328 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 111.395 0 112.515 1 ;
    END
  END Q[3]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.328 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 314.79 0 315.91 1 ;
    END
  END Q[4]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.328 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 355.545 0 356.665 1 ;
    END
  END Q[5]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.328 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 368.515 0 369.635 1 ;
    END
  END Q[6]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.328 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 409.275 0 410.395 1 ;
    END
  END Q[7]
  PIN WEN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
      ANTENNAGATEAREA 1.938 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 12.695 0 13.815 1 ;
    END
  END WEN[0]
  PIN WEN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
      ANTENNAGATEAREA 1.938 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 63.02 0 64.14 1 ;
    END
  END WEN[1]
  PIN WEN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
      ANTENNAGATEAREA 1.938 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 65.27 0 66.39 1 ;
    END
  END WEN[2]
  PIN WEN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
      ANTENNAGATEAREA 1.938 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 117.02 0 118.14 1 ;
    END
  END WEN[3]
  PIN WEN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
      ANTENNAGATEAREA 1.938 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 310.575 0 311.695 1 ;
    END
  END WEN[4]
  PIN WEN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
      ANTENNAGATEAREA 1.938 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 360.9 0 362.02 1 ;
    END
  END WEN[5]
  PIN WEN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
      ANTENNAGATEAREA 1.938 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 363.15 0 364.27 1 ;
    END
  END WEN[6]
  PIN WEN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
      ANTENNAGATEAREA 1.938 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 413.475 0 414.595 1 ;
    END
  END WEN[7]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 0 466.88 8.53 470.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 457.88 8.53 461.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 448.88 8.53 452.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 439.88 8.53 443.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 430.88 8.53 434.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 421.88 8.53 425.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 412.88 8.53 416.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 403.88 8.53 407.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 394.88 8.53 398.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 385.88 8.53 389.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 376.88 8.53 380.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 367.88 8.53 371.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 358.88 8.53 362.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 349.88 8.53 353.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 340.88 8.53 344.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 331.88 8.53 335.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 322.88 8.53 326.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 313.88 8.53 317.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 304.88 8.53 308.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 295.88 8.53 299.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 286.88 8.53 290.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 277.88 8.53 281.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 268.88 8.53 272.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 259.88 8.53 263.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 250.88 8.53 254.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 241.88 8.53 245.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 232.88 8.53 236.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 223.88 8.53 227.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 214.88 8.53 218.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 205.88 8.53 209.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 196.88 8.53 200.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 187.88 8.53 191.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 178.88 8.53 182.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 40.76 5.07 47.575 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 40.76 15.055 47.57 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 11.13 40.77 143.645 47.575 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 40.765 121.25 47.57 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 140.89 35.42 143.645 47.58 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 120.235 40.77 143.645 47.58 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 147.685 33.72 173.11 38.26 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 140.89 35.42 173.11 38.26 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 7.005 475.88 12.005 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 20.685 475.88 25.685 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 34.005 475.88 39.005 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 47.685 475.88 52.685 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 61.005 475.88 66.005 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.685 475.88 79.685 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 88.005 475.88 93.005 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 103.265 475.88 108.265 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 117.415 475.88 122.415 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 132.86 475.88 137.86 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 153.55 475.88 158.55 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 177.075 475.88 182.075 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 192.925 475.88 197.925 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 206.15 475.88 211.15 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 225.345 475.88 230.345 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 231.565 475.88 236.565 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 244.505 475.88 249.505 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 262.845 475.88 267.845 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 271.31 475.88 276.31 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 287.735 475.88 292.735 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 304.885 475.88 309.885 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 318.565 475.88 323.565 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 331.885 475.88 336.885 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 345.565 475.88 350.565 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 358.885 475.88 363.885 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 372.565 475.88 377.565 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 385.885 475.88 390.885 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 401.145 475.88 406.145 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 415.295 475.88 420.295 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 475.88 428.33 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 475.88 431.86 480.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 466.88 431.86 470.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 457.88 431.86 461.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 448.88 431.86 452.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 439.88 431.86 443.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 430.88 431.86 434.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 421.88 431.86 425.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 412.88 431.86 416.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 403.88 431.86 407.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 394.88 431.86 398.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 385.88 431.86 389.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 376.88 431.86 380.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 367.88 431.86 371.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 358.88 431.86 362.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 349.88 431.86 353.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 340.88 431.86 344.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 331.88 431.86 335.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 322.88 431.86 326.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 313.88 431.86 317.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 304.88 431.86 308.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 295.88 431.86 299.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 286.88 431.86 290.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 277.88 431.86 281.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 268.88 431.86 272.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 259.88 431.86 263.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 250.88 431.86 254.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 241.88 431.86 245.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 232.88 431.86 236.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 223.88 431.86 227.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 214.88 431.86 218.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 205.88 431.86 209.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 196.88 431.86 200.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 187.88 431.86 191.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 178.88 431.86 182.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 147.15 8.53 170.625 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 10.475 161.575 10.94 170.63 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 161.575 15.055 170.625 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 161.58 125.425 170.625 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 161.59 136.07 170.62 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 133.86 157.43 291.755 160.995 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 133.86 136.91 291.755 150.525 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 289.54 157.43 291.755 170.62 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 309.265 161.575 361.915 170.625 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 289.54 161.575 431.86 170.62 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 147.15 431.86 148.57 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 147.15 431.86 170.625 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 363.265 161.575 431.86 170.625 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 114.69 8.53 119.69 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 114.69 136.07 116.9 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 133.85 116.85 291.74 121.39 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 289.54 114.685 418.815 116.9 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 289.54 114.69 431.86 116.9 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 114.69 431.86 119.69 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 90.08 121.25 103.695 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 147.565 99.845 278.225 108.125 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 147.605 99.845 278.225 108.535 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 222.16 99.845 278.225 108.54 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 309.125 90.075 418.815 103.695 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 309.035 90.08 431.86 103.695 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 99.845 431.86 103.695 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 60.18 8.53 70.89 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 119.105 60.23 173.805 64.235 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 67.305 136.07 70.89 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 60.18 121.25 64.23 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 120.235 60.23 136.07 70.895 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 120.235 60.23 173.805 64.67 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 173.705 49.86 207.58 62.85 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 147.39 53.78 207.58 62.85 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 147.39 58.485 291.755 62.85 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 133.86 59.22 291.755 62.85 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 251.14 60.175 292.105 69.33 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 299.13 60.175 300.13 70.085 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 251.14 67.305 431.86 69.33 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 309.035 67.305 362.145 70.89 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 308.865 67.305 431.86 70.885 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 415.845 60.175 421.105 64.235 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 415.845 67.305 421.105 70.895 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 251.14 60.18 431.86 64.23 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 133.86 60.175 424.995 62.85 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 60.18 431.86 70.89 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 363.035 67.305 431.86 70.89 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 309.01 40.765 431.86 47.57 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 289.545 40.77 311.39 47.58 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 289.545 40.77 362.17 47.575 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 363.01 40.76 416.17 47.575 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 309.125 40.76 431.86 47.57 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 40.76 431.86 47.575 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 20.3 8.56 28.145 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 25.865 15.055 28.145 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 25.87 121.25 28.145 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 20.3 121.705 22.575 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 118.435 25.875 136.07 28.15 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 119.545 20.83 312.145 23.095 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 20.82 296.615 22.575 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 289.545 20.83 312.145 23.105 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 289.545 25.875 312.145 28.15 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 308.94 20.3 431.86 22.575 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 416.805 25.865 431.86 28.145 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 309.01 25.87 431.86 28.145 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.3 20.3 431.86 28.145 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 3.53 0 8.53 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 10.195 0 15.195 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 17.21 0 22.21 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 29.21 0 34.21 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 35.21 0 40.21 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 41.21 0 46.21 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 53.21 0 58.21 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 62.215 0 67.215 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 71.21 0 76.21 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 83.21 0 88.21 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 89.21 0 94.21 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 95.21 0 100.21 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 109.55 0 114.55 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 115.55 0 120.55 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 122.05 0 127.05 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 128.55 0 133.55 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 135.05 0 140.05 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 141.55 0 146.55 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 148.05 0 153.05 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 180.155 0 185.155 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 196.14 0 201.14 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 212.165 0 217.165 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 224.165 0 229.165 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 236.165 0 241.165 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 242.83 0 247.83 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 249.38 0 254.38 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 272.29 0 277.29 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 278.79 0 283.79 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 285.29 0 290.29 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 291.79 0 296.79 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 298.29 0 303.29 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 304.79 0 309.79 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 311.475 0 316.475 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 327.09 0 332.09 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 333.09 0 338.09 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 339.09 0 344.09 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 351.09 0 356.09 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 360.085 0 365.085 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 369.09 0 374.09 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 381.09 0 386.09 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 387.09 0 392.09 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 393.09 0 398.09 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 405.09 0 410.09 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 412.095 0 417.095 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 423.33 0 428.33 11.16 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 6.16 431.86 11.16 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 13.13 481.84 18.13 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 23.21 0 28.21 4.66 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 26.81 481.84 31.81 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 40.13 481.84 45.13 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 47.21 0 52.21 4.66 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 53.81 481.84 58.81 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 67.13 481.84 72.13 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 77.21 0 82.21 4.66 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 80.81 481.84 85.81 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 94.13 481.84 99.13 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 101.21 0 106.21 4.66 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 111.29 481.84 116.29 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 125.79 481.84 130.79 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 132.175 15.055 142.08 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 34.605 132.17 40.815 142.06 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 88.605 132.17 94.815 142.06 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 132.175 130.35 142.06 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 117.125 132.17 139.14 134.45 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 50.88 15.055 57.465 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 11.245 50.87 121.25 57.455 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 11.145 50.875 121.25 57.455 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 120.235 50.88 139.14 57.465 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 172.68 5.07 176.63 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 175.63 124.585 176.63 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 172.68 139.15 175.08 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 139.385 481.84 144.385 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 146.365 481.84 151.365 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 156.62 0 161.62 4.66 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 161.905 481.84 166.905 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 165.11 0 170.11 4.66 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 170.12 481.84 175.12 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 174.155 0 179.155 4.66 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 184.74 481.84 189.74 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 190.14 0 195.14 4.66 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 199.41 481.84 204.41 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 206.165 0 211.165 4.66 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 212.15 481.84 217.15 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 218.165 0 223.165 4.66 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 218.565 481.84 223.565 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 230.165 0 235.165 4.66 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 237.69 481.84 242.69 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 252.325 481.84 257.325 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 256.165 0 261.165 4.66 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 262.39 0 267.39 4.66 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 279.95 481.84 284.95 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 293.955 481.84 298.955 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 311.01 481.84 316.01 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 321.09 0 326.09 4.66 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 324.69 481.84 329.69 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 338.01 481.84 343.01 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 345.09 0 350.09 4.66 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 351.69 481.84 356.69 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 365.01 481.84 370.01 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 375.09 0 380.09 4.66 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 378.69 481.84 383.69 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 392.01 481.84 397.01 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 399.09 0 404.09 4.66 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 409.17 481.84 414.17 484.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 471.38 5.07 474.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 126.88 472.305 129.74 473.925 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 472.38 136.36 473.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.01 472.63 273.11 473.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 472.635 431.86 473.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 294.275 472.305 297.135 473.925 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 294.275 472.38 431.86 473.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 471.38 431.86 474.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 462.38 5.07 465.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 463.38 136.36 464.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 463.63 273.11 464.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 463.635 431.86 464.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 463.38 431.86 464.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 462.38 431.86 465.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 453.38 5.07 456.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 454.38 136.36 455.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 454.63 273.11 455.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 454.635 431.86 455.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 454.38 431.86 455.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 453.38 431.86 456.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 444.38 5.07 447.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 445.38 136.36 446.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 445.63 273.11 446.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 445.635 431.86 446.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 445.38 431.86 446.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 444.38 431.86 447.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 435.38 5.07 438.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 436.38 136.36 437.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 436.63 273.11 437.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 436.635 431.86 437.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 436.38 431.86 437.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 435.38 431.86 438.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 426.38 5.07 429.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 427.38 136.36 428.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 427.63 273.11 428.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 427.635 431.86 428.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 427.38 431.86 428.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 426.38 431.86 429.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 417.38 5.07 420.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 418.38 136.36 419.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 418.63 273.11 419.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 418.635 431.86 419.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 418.38 431.86 419.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 417.38 431.86 420.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 408.38 5.07 411.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 409.38 136.36 410.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 409.63 273.11 410.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 409.635 431.86 410.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 409.38 431.86 410.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 408.38 431.86 411.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 399.38 5.07 402.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 400.38 136.36 401.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 400.63 273.11 401.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 400.635 431.86 401.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 400.38 431.86 401.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 399.38 431.86 402.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 390.38 5.07 393.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 391.38 136.36 392.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 391.63 273.11 392.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 391.635 431.86 392.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 391.38 431.86 392.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 390.38 431.86 393.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 381.38 5.07 384.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 382.38 136.36 383.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 382.63 273.11 383.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 382.635 431.86 383.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 382.38 431.86 383.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 381.38 431.86 384.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 372.38 5.07 375.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 373.38 136.36 374.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 373.63 273.11 374.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 373.635 431.86 374.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 373.38 431.86 374.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 372.38 431.86 375.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 363.38 5.07 366.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 364.38 136.36 365.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 364.63 273.11 365.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 364.635 431.86 365.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 364.38 431.86 365.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 363.38 431.86 366.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 354.38 5.07 357.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 355.38 136.36 356.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 355.63 273.11 356.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 355.635 431.86 356.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 355.38 431.86 356.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 354.38 431.86 357.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 345.38 5.07 348.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 346.38 136.36 347.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 346.63 273.11 347.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 346.635 431.86 347.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 346.38 431.86 347.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 345.38 431.86 348.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 336.38 5.07 339.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 337.38 136.36 338.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 337.63 273.11 338.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 337.635 431.86 338.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 337.38 431.86 338.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 336.38 431.86 339.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 327.38 5.07 330.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 328.38 136.36 329.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 328.63 273.11 329.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 328.635 431.86 329.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 328.38 431.86 329.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 327.38 431.86 330.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 318.38 5.07 321.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 319.38 136.36 320.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 319.63 273.11 320.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 319.635 431.86 320.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 319.38 431.86 320.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 318.38 431.86 321.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 309.38 5.07 312.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 310.38 136.36 311.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 310.63 273.11 311.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 310.635 431.86 311.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 310.38 431.86 311.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 309.38 431.86 312.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 300.38 5.07 303.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 301.38 136.36 302.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 301.63 273.11 302.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 301.635 431.86 302.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 301.38 431.86 302.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 300.38 431.86 303.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 291.38 5.07 294.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 292.38 136.36 293.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 292.63 273.11 293.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 292.635 431.86 293.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 292.38 431.86 293.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 291.38 431.86 294.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 282.38 5.07 285.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 283.38 136.36 284.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 283.63 273.11 284.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 283.635 431.86 284.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 283.38 431.86 284.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 282.38 431.86 285.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 273.38 5.07 276.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 274.38 136.36 275.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 274.63 273.11 275.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 274.635 431.86 275.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 274.38 431.86 275.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 273.38 431.86 276.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 264.38 5.07 267.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 265.38 136.36 266.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 265.63 273.11 266.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 265.635 431.86 266.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 265.38 431.86 266.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 264.38 431.86 267.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 255.38 5.07 258.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 256.38 136.36 257.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 256.63 273.11 257.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 256.635 431.86 257.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 256.38 431.86 257.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 255.38 431.86 258.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 246.38 5.07 249.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 247.38 136.36 248.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 247.63 273.11 248.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 247.635 431.86 248.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 247.38 431.86 248.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 246.38 431.86 249.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 237.38 5.07 240.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 238.38 136.36 239.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 238.63 273.11 239.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 238.635 431.86 239.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 238.38 431.86 239.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 237.38 431.86 240.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 228.38 5.07 231.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 229.38 136.36 230.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 229.63 273.11 230.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 229.635 431.86 230.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 229.38 431.86 230.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 228.38 431.86 231.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 219.38 5.07 222.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 220.38 136.36 221.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 220.63 273.11 221.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 220.635 431.86 221.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 220.38 431.86 221.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 219.38 431.86 222.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 210.38 5.07 213.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 211.38 136.36 212.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 211.63 273.11 212.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 211.635 431.86 212.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 211.38 431.86 212.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 210.38 431.86 213.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 201.38 5.07 204.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 202.38 136.36 203.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 202.63 273.11 203.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 202.635 431.86 203.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 202.38 431.86 203.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 201.38 431.86 204.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 192.38 5.07 195.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 193.38 136.36 194.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 193.63 273.11 194.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 193.635 431.86 194.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 193.38 431.86 194.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 192.38 431.86 195.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 183.38 5.07 186.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 184.38 136.36 185.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 184.63 273.11 185.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 184.635 431.86 185.64 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.105 184.38 431.86 185.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 183.38 431.86 186.88 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 302.3 175.79 431.86 176.49 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 293.955 172.68 431.86 175.08 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 172.68 431.86 176.63 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 416.8 175.63 431.86 176.63 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 286.475 132.175 431.86 134.45 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 332.485 132.17 338.695 142.06 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 386.485 132.17 392.695 142.06 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 293.925 132.175 431.86 142.06 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 416.805 132.175 431.86 142.08 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 106.41 5.07 111.41 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 120.18 109.13 139.13 111.41 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 109.135 139.13 111.41 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 136.935 109.13 139.13 115.995 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 280.39 109.13 288.405 115.995 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 136.935 111.455 288.405 115.995 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 280.39 109.13 418.815 111.41 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 106.41 431.86 111.41 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 280.39 109.135 431.86 111.41 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 71.64 118.39 88.65 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 71.64 121.25 82.985 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 120.555 71.645 139.14 82.99 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 147.39 66.215 229.885 75.075 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 136.935 66.225 229.885 75.075 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 72.455 238.415 75.075 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 207.465 65.39 248.875 68.8 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 74.68 258.8 75.075 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 74.83 278.225 75.075 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 234.91 74.84 431.86 83.92 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 286.475 71.635 418.815 83.92 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 309.035 71.64 431.86 88.65 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 286.475 50.88 431.86 57.455 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 211.305 53.7 431.86 57.455 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 309.125 50.865 422.41 57.465 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 309.025 50.875 422.41 57.455 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 309.125 50.88 431.86 57.465 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 28.83 5.07 37.98 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 28.83 15.055 30.995 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 34.91 15.055 37.98 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 11.245 34.9 121.25 37.975 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 11.13 34.905 121.25 37.975 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 118.125 34.91 139.14 37.98 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 118.435 30.885 206.985 30.995 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 147.29 28.325 173.11 32.865 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 28.83 173.11 30.99 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 147.29 30.885 206.985 32.865 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 174.3 30.885 206.985 42.91 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 147.565 39.5 206.985 42.91 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 174.3 32.96 277.41 36.96 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 209.285 45.825 257.15 52.1 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 254.61 28.025 277.41 47.51 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 254.61 34.92 288.68 44.65 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 254.61 28.83 312.145 30.995 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 254.61 34.92 313.735 37.98 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 254.61 28.83 431.86 30.99 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 309.125 34.9 423.935 37.975 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 309.01 34.905 423.935 37.975 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 416.805 28.83 431.86 30.995 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 28.83 431.86 37.98 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 416.805 34.91 431.86 37.98 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 12.51 5.07 18.86 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 17.1 15.055 18.86 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 17.105 121.705 18.86 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 137.19 17.62 138.89 19.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 143.82 17.62 144.47 19.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 208.87 17.62 209.52 19.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 211.495 17.62 212.145 19.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 234.365 17.62 235.015 19.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 236.605 17.62 237.255 19.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 238.845 17.62 239.495 19.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 241.085 17.62 241.735 19.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 119.545 17.62 306.075 19.375 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 286.725 17.62 306.075 19.38 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 12.51 431.86 14.27 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 304.43 17.1 431.86 18.86 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 426.79 12.51 431.86 18.86 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0 0 431.86 484.88 ;
    LAYER Metal2 ;
      POLYGON 431.86 484.88 0 484.88 0 0 9.04 0 9.04 1.28 10.72 1.28 10.72 0 12.415 0 12.415 1.28 14.095 1.28 14.095 0 16.62 0 16.62 1.28 18.3 1.28 18.3 0 57.385 0 57.385 1.28 59.065 1.28 59.065 0 60.75 0 60.75 1.28 62.43 1.28 62.43 0 62.74 0 62.74 1.28 64.42 1.28 64.42 0 64.99 0 64.99 1.28 66.67 1.28 66.67 0 66.99 0 66.99 1.28 68.67 1.28 68.67 0 70.355 0 70.355 1.28 72.035 1.28 72.035 0 111.115 0 111.115 1.28 112.795 1.28 112.795 0 116.74 0 116.74 1.28 118.42 1.28 118.42 0 118.695 0 118.695 1.28 120.375 1.28 120.375 0 139.4 0 139.4 1.28 141.08 1.28 141.08 0 144.75 0 144.75 1.28 146.43 1.28 146.43 0 148.245 0 148.245 1.28 149.925 1.28 149.925 0 154.015 0 154.015 1.28 155.695 1.28 155.695 0 162.48 0 162.48 1.28 164.16 1.28 164.16 0 170.935 0 170.935 1.28 172.615 1.28 172.615 0 202.66 0 202.66 1.28 204.34 1.28 204.34 0 251.43 0 251.43 1.28 253.11 1.28 253.11 0 268.58 0 268.58 1.28 270.26 1.28 270.26 0 271.805 0 271.805 1.28 273.485 1.28 273.485 0 275.54 0 275.54 1.28 277.22 1.28 277.22 0 281.045 0 281.045 1.28 282.725 1.28 282.725 0 306.955 0 306.955 1.28 308.635 1.28 308.635 0 310.295 0 310.295 1.28 311.975 1.28 311.975 0 314.51 0 314.51 1.28 316.19 1.28 316.19 0 355.265 0 355.265 1.28 356.945 1.28 356.945 0 358.63 0 358.63 1.28 360.31 1.28 360.31 0 360.62 0 360.62 1.28 362.3 1.28 362.3 0 362.87 0 362.87 1.28 364.55 1.28 364.55 0 364.87 0 364.87 1.28 366.55 1.28 366.55 0 368.235 0 368.235 1.28 369.915 1.28 369.915 0 408.995 0 408.995 1.28 410.675 1.28 410.675 0 413.195 0 413.195 1.28 414.875 1.28 414.875 0 416.58 0 416.58 1.28 418.26 1.28 418.26 0 431.86 0 ;
    LAYER Via1 ;
      RECT 0 0 431.86 484.88 ;
    LAYER Via2 ;
      RECT 0 0 431.86 484.88 ;
    LAYER Metal3 ;
      POLYGON 400.865 484.88 397.29 484.88 397.29 481.56 391.73 481.56 391.73 484.88 391.165 484.88 391.165 481.16 400.865 481.16 ;
      RECT 356.37 0 359.805 5.88 ;
      RECT 127.33 0 128.27 5.88 ;
      POLYGON 431.86 89.8 419.095 89.8 419.095 89.795 308.845 89.795 308.845 89.8 308.755 89.8 308.755 99.565 121.53 99.565 121.53 89.8 0 89.8 0 88.93 118.67 88.93 118.67 83.265 120.275 83.265 120.275 83.27 139.42 83.27 139.42 75.355 234.63 75.355 234.63 84.2 308.755 84.2 308.755 88.93 431.86 88.93 ;
      RECT 417.375 0 423.05 5.88 ;
      POLYGON 431.86 214.6 423.05 214.6 423.05 218.66 431.86 218.66 431.86 219.1 426.51 219.1 426.51 220.1 296.825 220.1 296.825 220.355 273.39 220.355 273.39 220.35 151.735 220.35 151.735 220.355 136.64 220.355 136.64 220.1 5.35 220.1 5.35 219.1 0 219.1 0 218.66 8.81 218.66 8.81 214.6 0 214.6 0 214.16 5.35 214.16 5.35 213.16 136.64 213.16 136.64 212.92 296.825 212.92 296.825 213.16 426.51 213.16 426.51 214.16 431.86 214.16 ;
      RECT 230.625 481.16 231.285 484.88 ;
      RECT 338.37 0 338.81 5.88 ;
      RECT 114.83 0 115.27 5.88 ;
      POLYGON 431.86 286.6 423.05 286.6 423.05 290.66 431.86 290.66 431.86 291.1 426.51 291.1 426.51 292.1 296.825 292.1 296.825 292.355 273.39 292.355 273.39 292.35 151.735 292.35 151.735 292.355 136.64 292.355 136.64 292.1 5.35 292.1 5.35 291.1 0 291.1 0 290.66 8.81 290.66 8.81 286.6 0 286.6 0 286.16 5.35 286.16 5.35 285.16 136.64 285.16 136.64 284.92 296.825 284.92 296.825 285.16 426.51 285.16 426.51 286.16 431.86 286.16 ;
      POLYGON 423.05 67.025 300.41 67.025 300.41 64.51 415.565 64.51 415.565 64.515 421.385 64.515 421.385 64.51 423.05 64.51 ;
      RECT 290.57 0 291.51 5.88 ;
      POLYGON 223.885 5.88 217.445 5.88 217.445 0 217.885 0 217.885 4.94 223.445 4.94 223.445 0 223.885 0 ;
      POLYGON 385.605 484.88 383.97 484.88 383.97 481.56 378.41 481.56 378.41 484.88 377.845 484.88 377.845 481.16 385.605 481.16 ;
      POLYGON 431.86 304.6 423.05 304.6 423.05 308.66 431.86 308.66 431.86 309.1 426.51 309.1 426.51 310.1 296.825 310.1 296.825 310.355 273.39 310.355 273.39 310.35 151.735 310.35 151.735 310.355 136.64 310.355 136.64 310.1 5.35 310.1 5.35 309.1 0 309.1 0 308.66 8.81 308.66 8.81 304.6 0 304.6 0 304.16 5.35 304.16 5.35 303.16 136.64 303.16 136.64 302.92 296.825 302.92 296.825 303.16 426.51 303.16 426.51 304.16 431.86 304.16 ;
      POLYGON 431.86 131.895 392.975 131.895 392.975 131.89 386.205 131.89 386.205 131.895 338.975 131.895 338.975 131.89 332.205 131.89 332.205 131.895 286.195 131.895 286.195 134.73 293.645 134.73 293.645 142.34 416.525 142.34 416.525 142.36 431.86 142.36 431.86 146.87 292.035 146.87 292.035 136.63 133.58 136.63 133.58 146.87 0 146.87 0 142.36 15.335 142.36 15.335 142.34 130.63 142.34 130.63 134.73 139.42 134.73 139.42 131.89 116.845 131.89 116.845 131.895 95.095 131.895 95.095 131.89 88.325 131.89 88.325 131.895 41.095 131.895 41.095 131.89 34.325 131.89 34.325 131.895 0 131.895 0 119.97 8.81 119.97 8.81 117.18 133.57 117.18 133.57 121.67 292.02 121.67 292.02 117.18 423.05 117.18 423.05 119.97 431.86 119.97 ;
      POLYGON 431.86 439.6 423.05 439.6 423.05 443.66 431.86 443.66 431.86 444.1 426.51 444.1 426.51 445.1 296.825 445.1 296.825 445.355 273.39 445.355 273.39 445.35 151.735 445.35 151.735 445.355 136.64 445.355 136.64 445.1 5.35 445.1 5.35 444.1 0 444.1 0 443.66 8.81 443.66 8.81 439.6 0 439.6 0 439.16 5.35 439.16 5.35 438.16 136.64 438.16 136.64 437.92 296.825 437.92 296.825 438.16 426.51 438.16 426.51 439.16 431.86 439.16 ;
      POLYGON 431.86 295.6 423.05 295.6 423.05 299.66 431.86 299.66 431.86 300.1 426.51 300.1 426.51 301.1 296.825 301.1 296.825 301.355 273.39 301.355 273.39 301.35 151.735 301.35 151.735 301.355 136.64 301.355 136.64 301.1 5.35 301.1 5.35 300.1 0 300.1 0 299.66 8.81 299.66 8.81 295.6 0 295.6 0 295.16 5.35 295.16 5.35 294.16 136.64 294.16 136.64 293.92 296.825 293.92 296.825 294.16 426.51 294.16 426.51 295.16 431.86 295.16 ;
      RECT 0 0 3.25 5.88 ;
      RECT 34.49 0 34.93 5.88 ;
      POLYGON 225.065 484.88 223.845 484.88 223.845 481.56 218.285 481.56 218.285 484.88 217.43 484.88 217.43 481.56 211.87 481.56 211.87 484.88 211.43 484.88 211.43 481.16 225.065 481.16 ;
      RECT 0 481.16 6.725 484.88 ;
      POLYGON 153.27 484.88 151.645 484.88 151.645 481.56 146.085 481.56 146.085 484.88 144.665 484.88 144.665 481.56 139.105 481.56 139.105 484.88 138.14 484.88 138.14 481.16 153.27 481.16 ;
      POLYGON 431.86 331.6 423.05 331.6 423.05 335.66 431.86 335.66 431.86 336.1 426.51 336.1 426.51 337.1 296.825 337.1 296.825 337.355 273.39 337.355 273.39 337.35 151.735 337.35 151.735 337.355 136.64 337.355 136.64 337.1 5.35 337.1 5.35 336.1 0 336.1 0 335.66 8.81 335.66 8.81 331.6 0 331.6 0 331.16 5.35 331.16 5.35 330.16 136.64 330.16 136.64 329.92 296.825 329.92 296.825 330.16 426.51 330.16 426.51 331.16 431.86 331.16 ;
      POLYGON 404.81 5.88 398.37 5.88 398.37 0 398.81 0 398.81 4.94 404.37 4.94 404.37 0 404.81 0 ;
      RECT 284.07 0 285.01 5.88 ;
      RECT 88.49 0 88.93 5.88 ;
      POLYGON 272.01 5.88 254.66 5.88 254.66 0 255.885 0 255.885 4.94 261.445 4.94 261.445 0 262.11 0 262.11 4.94 267.67 4.94 267.67 0 272.01 0 ;
      POLYGON 211.885 5.88 201.42 5.88 201.42 0 205.885 0 205.885 4.94 211.445 4.94 211.445 0 211.885 0 ;
      POLYGON 372.285 484.88 370.29 484.88 370.29 481.56 364.73 481.56 364.73 484.88 364.165 484.88 364.165 481.16 372.285 481.16 ;
      POLYGON 431.86 223.6 423.05 223.6 423.05 227.66 431.86 227.66 431.86 228.1 426.51 228.1 426.51 229.1 296.825 229.1 296.825 229.355 273.39 229.355 273.39 229.35 151.735 229.35 151.735 229.355 136.64 229.355 136.64 229.1 5.35 229.1 5.35 228.1 0 228.1 0 227.66 8.81 227.66 8.81 223.6 0 223.6 0 223.16 5.35 223.16 5.35 222.16 136.64 222.16 136.64 221.92 296.825 221.92 296.825 222.16 426.51 222.16 426.51 223.16 431.86 223.16 ;
      RECT 140.33 0 141.27 5.88 ;
      POLYGON 179.875 5.88 153.33 5.88 153.33 0 156.34 0 156.34 4.94 161.9 4.94 161.9 0 164.83 0 164.83 4.94 170.39 4.94 170.39 0 173.875 0 173.875 4.94 179.435 4.94 179.435 0 179.875 0 ;
      POLYGON 431.86 232.6 423.05 232.6 423.05 236.66 431.86 236.66 431.86 237.1 426.51 237.1 426.51 238.1 296.825 238.1 296.825 238.355 273.39 238.355 273.39 238.35 151.735 238.35 151.735 238.355 136.64 238.355 136.64 238.1 5.35 238.1 5.35 237.1 0 237.1 0 236.66 8.81 236.66 8.81 232.6 0 232.6 0 232.16 5.35 232.16 5.35 231.16 136.64 231.16 136.64 230.92 296.825 230.92 296.825 231.16 426.51 231.16 426.51 232.16 431.86 232.16 ;
      POLYGON 431.86 421.6 423.05 421.6 423.05 425.66 431.86 425.66 431.86 426.1 426.51 426.1 426.51 427.1 296.825 427.1 296.825 427.355 273.39 427.355 273.39 427.35 151.735 427.35 151.735 427.355 136.64 427.355 136.64 427.1 5.35 427.1 5.35 426.1 0 426.1 0 425.66 8.81 425.66 8.81 421.6 0 421.6 0 421.16 5.35 421.16 5.35 420.16 136.64 420.16 136.64 419.92 296.825 419.92 296.825 420.16 426.51 420.16 426.51 421.16 431.86 421.16 ;
      POLYGON 87.725 484.88 86.09 484.88 86.09 481.56 80.53 481.56 80.53 484.88 79.965 484.88 79.965 481.16 87.725 481.16 ;
      POLYGON 431.86 250.6 423.05 250.6 423.05 254.66 431.86 254.66 431.86 255.1 426.51 255.1 426.51 256.1 296.825 256.1 296.825 256.355 273.39 256.355 273.39 256.35 151.735 256.35 151.735 256.355 136.64 256.355 136.64 256.1 5.35 256.1 5.35 255.1 0 255.1 0 254.66 8.81 254.66 8.81 250.6 0 250.6 0 250.16 5.35 250.16 5.35 249.16 136.64 249.16 136.64 248.92 296.825 248.92 296.825 249.16 426.51 249.16 426.51 250.16 431.86 250.16 ;
      RECT 0 11.44 431.86 12.23 ;
      POLYGON 119.955 67.025 8.81 67.025 8.81 64.51 118.825 64.51 118.825 64.515 119.955 64.515 ;
      RECT 303.57 0 304.51 5.88 ;
      POLYGON 74.405 484.88 72.41 484.88 72.41 481.56 66.85 481.56 66.85 484.88 66.285 484.88 66.285 481.16 74.405 481.16 ;
      RECT 428.61 481.16 431.86 484.88 ;
      RECT 297.07 0 298.01 5.88 ;
      RECT 420.575 481.16 423.05 484.88 ;
      POLYGON 20.405 484.88 18.41 484.88 18.41 481.56 12.85 481.56 12.85 484.88 12.285 484.88 12.285 481.16 20.405 481.16 ;
      POLYGON 304.605 484.88 299.235 484.88 299.235 481.56 293.675 481.56 293.675 484.88 293.015 484.88 293.015 481.16 304.605 481.16 ;
      POLYGON 431.86 187.6 423.05 187.6 423.05 191.66 431.86 191.66 431.86 192.1 426.51 192.1 426.51 193.1 296.825 193.1 296.825 193.355 273.39 193.355 273.39 193.35 151.735 193.35 151.735 193.355 136.64 193.355 136.64 193.1 5.35 193.1 5.35 192.1 0 192.1 0 191.66 8.81 191.66 8.81 187.6 0 187.6 0 187.16 5.35 187.16 5.35 186.16 136.64 186.16 136.64 185.92 296.825 185.92 296.825 186.16 426.51 186.16 426.51 187.16 431.86 187.16 ;
      POLYGON 431.86 196.6 423.05 196.6 423.05 200.66 431.86 200.66 431.86 201.1 426.51 201.1 426.51 202.1 296.825 202.1 296.825 202.355 273.39 202.355 273.39 202.35 151.735 202.35 151.735 202.355 136.64 202.355 136.64 202.1 5.35 202.1 5.35 201.1 0 201.1 0 200.66 8.81 200.66 8.81 196.6 0 196.6 0 196.16 5.35 196.16 5.35 195.16 136.64 195.16 136.64 194.92 296.825 194.92 296.825 195.16 426.51 195.16 426.51 196.16 431.86 196.16 ;
      RECT 58.49 0 61.935 5.88 ;
      POLYGON 318.285 484.88 316.29 484.88 316.29 481.56 310.73 481.56 310.73 484.88 310.165 484.88 310.165 481.16 318.285 481.16 ;
      RECT 248.11 0 249.1 5.88 ;
      POLYGON 358.605 484.88 356.97 484.88 356.97 481.56 351.41 481.56 351.41 484.88 350.845 484.88 350.845 481.16 358.605 481.16 ;
      POLYGON 431.86 241.6 423.05 241.6 423.05 245.66 431.86 245.66 431.86 246.1 426.51 246.1 426.51 247.1 296.825 247.1 296.825 247.355 273.39 247.355 273.39 247.35 151.735 247.35 151.735 247.355 136.64 247.355 136.64 247.1 5.35 247.1 5.35 246.1 0 246.1 0 245.66 8.81 245.66 8.81 241.6 0 241.6 0 241.16 5.35 241.16 5.35 240.16 136.64 240.16 136.64 239.92 296.825 239.92 296.825 240.16 426.51 240.16 426.51 241.16 431.86 241.16 ;
      POLYGON 60.725 484.88 59.09 484.88 59.09 481.56 53.53 481.56 53.53 484.88 52.965 484.88 52.965 481.16 60.725 481.16 ;
      POLYGON 82.93 5.88 76.49 5.88 76.49 0 76.93 0 76.93 4.94 82.49 4.94 82.49 0 82.93 0 ;
      POLYGON 350.81 5.88 344.37 5.88 344.37 0 344.81 0 344.81 4.94 350.37 4.94 350.37 0 350.81 0 ;
      POLYGON 47.405 484.88 45.41 484.88 45.41 481.56 39.85 481.56 39.85 484.88 39.285 484.88 39.285 481.16 47.405 481.16 ;
      POLYGON 431.86 466.6 423.05 466.6 423.05 470.66 431.86 470.66 431.86 471.1 426.51 471.1 426.51 472.1 297.415 472.1 297.415 472.025 293.995 472.025 293.995 472.355 273.39 472.355 273.39 472.35 151.73 472.35 151.73 472.355 136.64 472.355 136.64 472.1 130.02 472.1 130.02 472.025 126.6 472.025 126.6 472.1 5.35 472.1 5.35 471.1 0 471.1 0 470.66 8.81 470.66 8.81 466.6 0 466.6 0 466.16 5.35 466.16 5.35 465.16 136.64 465.16 136.64 464.92 296.825 464.92 296.825 465.16 426.51 465.16 426.51 466.16 431.86 466.16 ;
      POLYGON 132.58 484.88 131.07 484.88 131.07 481.56 125.51 481.56 125.51 484.88 122.695 484.88 122.695 481.16 132.58 481.16 ;
      POLYGON 431.86 172.4 293.675 172.4 293.675 175.36 416.52 175.36 416.52 175.51 302.02 175.51 302.02 176.77 416.52 176.77 416.52 176.91 431.86 176.91 431.86 178.6 423.05 178.6 423.05 182.66 431.86 182.66 431.86 183.1 426.51 183.1 426.51 184.1 296.825 184.1 296.825 184.355 273.39 184.355 273.39 184.35 151.735 184.35 151.735 184.355 136.64 184.355 136.64 184.1 5.35 184.1 5.35 183.1 0 183.1 0 182.66 8.81 182.66 8.81 178.6 0 178.6 0 176.91 124.865 176.91 124.865 175.36 139.43 175.36 139.43 172.4 0 172.4 0 170.905 10.195 170.905 10.195 170.91 11.22 170.91 11.22 170.905 125.705 170.905 125.705 170.9 136.35 170.9 136.35 161.31 125.705 161.31 125.705 161.3 15.335 161.3 15.335 161.295 8.81 161.295 8.81 148.85 133.58 148.85 133.58 150.805 292.035 150.805 292.035 148.85 423.05 148.85 423.05 161.295 292.035 161.295 292.035 157.15 133.58 157.15 133.58 161.275 289.26 161.275 289.26 170.9 308.985 170.9 308.985 170.905 362.195 170.905 362.195 170.9 362.985 170.9 362.985 170.905 431.86 170.905 ;
      POLYGON 109.27 5.88 100.49 5.88 100.49 0 100.93 0 100.93 4.94 106.49 4.94 106.49 0 109.27 0 ;
      RECT 120.83 0 121.77 5.88 ;
      RECT 133.83 0 134.77 5.88 ;
      POLYGON 431.86 205.6 423.05 205.6 423.05 209.66 431.86 209.66 431.86 210.1 426.51 210.1 426.51 211.1 296.825 211.1 296.825 211.355 273.39 211.355 273.39 211.35 151.735 211.35 151.735 211.355 136.64 211.355 136.64 211.1 5.35 211.1 5.35 210.1 0 210.1 0 209.66 8.81 209.66 8.81 205.6 0 205.6 0 205.16 5.35 205.16 5.35 204.16 136.64 204.16 136.64 203.92 296.825 203.92 296.825 204.16 426.51 204.16 426.51 205.16 431.86 205.16 ;
      RECT 94.49 0 94.93 5.88 ;
      RECT 392.37 0 392.81 5.88 ;
      POLYGON 380.81 5.88 374.37 5.88 374.37 0 374.81 0 374.81 4.94 380.37 4.94 380.37 0 380.81 0 ;
      POLYGON 102.985 484.88 99.41 484.88 99.41 481.56 93.85 481.56 93.85 484.88 93.285 484.88 93.285 481.16 102.985 481.16 ;
      RECT 365.365 0 368.81 5.88 ;
      POLYGON 431.86 313.6 423.05 313.6 423.05 317.66 431.86 317.66 431.86 318.1 426.51 318.1 426.51 319.1 296.825 319.1 296.825 319.355 273.39 319.355 273.39 319.35 151.735 319.35 151.735 319.355 136.64 319.355 136.64 319.1 5.35 319.1 5.35 318.1 0 318.1 0 317.66 8.81 317.66 8.81 313.6 0 313.6 0 313.16 5.35 313.16 5.35 312.16 136.64 312.16 136.64 311.92 296.825 311.92 296.825 312.16 426.51 312.16 426.51 313.16 431.86 313.16 ;
      POLYGON 326.81 5.88 316.755 5.88 316.755 0 320.81 0 320.81 4.94 326.37 4.94 326.37 0 326.81 0 ;
      POLYGON 431.86 322.6 423.05 322.6 423.05 326.66 431.86 326.66 431.86 327.1 426.51 327.1 426.51 328.1 296.825 328.1 296.825 328.355 273.39 328.355 273.39 328.35 151.735 328.35 151.735 328.355 136.64 328.355 136.64 328.1 5.35 328.1 5.35 327.1 0 327.1 0 326.66 8.81 326.66 8.81 322.6 0 322.6 0 322.16 5.35 322.16 5.35 321.16 136.64 321.16 136.64 320.92 296.825 320.92 296.825 321.16 426.51 321.16 426.51 322.16 431.86 322.16 ;
      POLYGON 431.86 114.41 419.095 114.41 419.095 114.405 289.26 114.405 289.26 116.57 136.35 116.57 136.35 114.41 0 114.41 0 111.69 136.655 111.69 136.655 116.275 288.685 116.275 288.685 111.69 431.86 111.69 ;
      RECT 40.49 0 40.93 5.88 ;
      POLYGON 235.885 5.88 229.445 5.88 229.445 0 229.885 0 229.885 4.94 235.445 4.94 235.445 0 235.885 0 ;
      POLYGON 431.86 367.6 423.05 367.6 423.05 371.66 431.86 371.66 431.86 372.1 426.51 372.1 426.51 373.1 296.825 373.1 296.825 373.355 273.39 373.355 273.39 373.35 151.735 373.35 151.735 373.355 136.64 373.355 136.64 373.1 5.35 373.1 5.35 372.1 0 372.1 0 371.66 8.81 371.66 8.81 367.6 0 367.6 0 367.16 5.35 367.16 5.35 366.16 136.64 366.16 136.64 365.92 296.825 365.92 296.825 366.16 426.51 366.16 426.51 367.16 431.86 367.16 ;
      POLYGON 331.605 484.88 329.97 484.88 329.97 481.56 324.41 481.56 324.41 484.88 323.845 484.88 323.845 481.16 331.605 481.16 ;
      RECT 268.125 481.16 271.03 484.88 ;
      POLYGON 192.645 484.88 190.02 484.88 190.02 481.56 184.46 481.56 184.46 484.88 182.355 484.88 182.355 481.16 192.645 481.16 ;
      RECT 292.385 64.51 298.85 67.025 ;
      POLYGON 28.93 5.88 22.49 5.88 22.49 0 22.93 0 22.93 4.94 28.49 4.94 28.49 0 28.93 0 ;
      POLYGON 205.87 484.88 204.69 484.88 204.69 481.56 199.13 481.56 199.13 484.88 198.205 484.88 198.205 481.16 205.87 481.16 ;
      POLYGON 431.86 430.6 423.05 430.6 423.05 434.66 431.86 434.66 431.86 435.1 426.51 435.1 426.51 436.1 296.825 436.1 296.825 436.355 273.39 436.355 273.39 436.35 151.735 436.35 151.735 436.355 136.64 436.355 136.64 436.1 5.35 436.1 5.35 435.1 0 435.1 0 434.66 8.81 434.66 8.81 430.6 0 430.6 0 430.16 5.35 430.16 5.35 429.16 136.64 429.16 136.64 428.92 296.825 428.92 296.825 429.16 426.51 429.16 426.51 430.16 431.86 430.16 ;
      POLYGON 52.93 5.88 46.49 5.88 46.49 0 46.93 0 46.93 4.94 52.49 4.94 52.49 0 52.93 0 ;
      POLYGON 415.015 484.88 414.45 484.88 414.45 481.56 408.89 481.56 408.89 484.88 406.425 484.88 406.425 481.16 415.015 481.16 ;
      POLYGON 431.86 358.6 423.05 358.6 423.05 362.66 431.86 362.66 431.86 363.1 426.51 363.1 426.51 364.1 296.825 364.1 296.825 364.355 273.39 364.355 273.39 364.35 151.735 364.35 151.735 364.355 136.64 364.355 136.64 364.1 5.35 364.1 5.35 363.1 0 363.1 0 362.66 8.81 362.66 8.81 358.6 0 358.6 0 358.16 5.35 358.16 5.35 357.16 136.64 357.16 136.64 356.92 296.825 356.92 296.825 357.16 426.51 357.16 426.51 358.16 431.86 358.16 ;
      POLYGON 431.86 457.6 423.05 457.6 423.05 461.66 431.86 461.66 431.86 462.1 426.51 462.1 426.51 463.1 296.825 463.1 296.825 463.355 273.39 463.355 273.39 463.35 151.735 463.35 151.735 463.355 136.64 463.355 136.64 463.1 5.35 463.1 5.35 462.1 0 462.1 0 461.66 8.81 461.66 8.81 457.6 0 457.6 0 457.16 5.35 457.16 5.35 456.16 136.64 456.16 136.64 455.92 296.825 455.92 296.825 456.16 426.51 456.16 426.51 457.16 431.86 457.16 ;
      POLYGON 431.86 340.6 423.05 340.6 423.05 344.66 431.86 344.66 431.86 345.1 426.51 345.1 426.51 346.1 296.825 346.1 296.825 346.355 273.39 346.355 273.39 346.35 151.735 346.35 151.735 346.355 136.64 346.355 136.64 346.1 5.35 346.1 5.35 345.1 0 345.1 0 344.66 8.81 344.66 8.81 340.6 0 340.6 0 340.16 5.35 340.16 5.35 339.16 136.64 339.16 136.64 338.92 296.825 338.92 296.825 339.16 426.51 339.16 426.51 340.16 431.86 340.16 ;
      POLYGON 431.86 349.6 423.05 349.6 423.05 353.66 431.86 353.66 431.86 354.1 426.51 354.1 426.51 355.1 296.825 355.1 296.825 355.355 273.39 355.355 273.39 355.35 151.735 355.35 151.735 355.355 136.64 355.355 136.64 355.1 5.35 355.1 5.35 354.1 0 354.1 0 353.66 8.81 353.66 8.81 349.6 0 349.6 0 349.16 5.35 349.16 5.35 348.16 136.64 348.16 136.64 347.92 296.825 347.92 296.825 348.16 426.51 348.16 426.51 349.16 431.86 349.16 ;
      RECT 332.37 0 332.81 5.88 ;
      POLYGON 262.565 484.88 257.605 484.88 257.605 481.56 252.045 481.56 252.045 484.88 249.785 484.88 249.785 481.16 262.565 481.16 ;
      RECT 15.475 0 16.93 5.88 ;
      RECT 67.495 0 70.93 5.88 ;
      POLYGON 431.86 20.02 308.66 20.02 308.66 20.55 296.895 20.55 296.895 20.54 121.985 20.54 121.985 20.02 0 20.02 0 19.14 119.265 19.14 119.265 19.655 136.91 19.655 136.91 19.66 139.17 19.66 139.17 19.655 143.54 19.655 143.54 19.66 144.75 19.66 144.75 19.655 208.59 19.655 208.59 19.66 209.8 19.66 209.8 19.655 211.215 19.655 211.215 19.66 212.425 19.66 212.425 19.655 234.085 19.655 234.085 19.66 235.295 19.66 235.295 19.655 236.325 19.655 236.325 19.66 237.535 19.66 237.535 19.655 238.565 19.655 238.565 19.66 239.775 19.66 239.775 19.655 240.805 19.655 240.805 19.66 242.015 19.66 242.015 19.655 286.445 19.655 286.445 19.66 306.355 19.66 306.355 19.14 431.86 19.14 ;
      RECT 146.83 0 147.77 5.88 ;
      POLYGON 431.86 71.36 419.095 71.36 419.095 71.355 286.195 71.355 286.195 74.56 278.505 74.56 278.505 74.55 259.08 74.55 259.08 74.4 238.695 74.4 238.695 72.175 230.165 72.175 230.165 69.08 249.155 69.08 249.155 65.11 207.185 65.11 207.185 65.935 147.11 65.935 147.11 65.945 136.655 65.945 136.655 71.365 121.53 71.365 121.53 71.36 0 71.36 0 71.17 119.955 71.17 119.955 71.175 136.35 71.175 136.35 64.95 174.085 64.95 174.085 63.13 250.86 63.13 250.86 69.61 298.85 69.61 298.85 70.365 300.41 70.365 300.41 69.61 308.585 69.61 308.585 71.165 308.755 71.165 308.755 71.17 362.425 71.17 362.425 71.165 362.755 71.165 362.755 71.17 415.565 71.17 415.565 71.175 421.385 71.175 421.385 71.17 431.86 71.17 ;
      POLYGON 426.51 16.82 304.15 16.82 304.15 17.34 121.985 17.34 121.985 16.825 15.335 16.825 15.335 16.82 5.35 16.82 5.35 14.55 426.51 14.55 ;
      RECT 428.61 0 431.86 5.88 ;
      POLYGON 431.86 448.6 423.05 448.6 423.05 452.66 431.86 452.66 431.86 453.1 426.51 453.1 426.51 454.1 296.825 454.1 296.825 454.355 273.39 454.355 273.39 454.35 151.735 454.35 151.735 454.355 136.64 454.355 136.64 454.1 5.35 454.1 5.35 453.1 0 453.1 0 452.66 8.81 452.66 8.81 448.6 0 448.6 0 448.16 5.35 448.16 5.35 447.16 136.64 447.16 136.64 446.92 296.825 446.92 296.825 447.16 426.51 447.16 426.51 448.16 431.86 448.16 ;
      RECT 8.81 0 9.915 5.88 ;
      POLYGON 431.86 394.6 423.05 394.6 423.05 398.66 431.86 398.66 431.86 399.1 426.51 399.1 426.51 400.1 296.825 400.1 296.825 400.355 273.39 400.355 273.39 400.35 151.735 400.35 151.735 400.355 136.64 400.355 136.64 400.1 5.35 400.1 5.35 399.1 0 399.1 0 398.66 8.81 398.66 8.81 394.6 0 394.6 0 394.16 5.35 394.16 5.35 393.16 136.64 393.16 136.64 392.92 296.825 392.92 296.825 393.16 426.51 393.16 426.51 394.16 431.86 394.16 ;
      POLYGON 431.86 412.6 423.05 412.6 423.05 416.66 431.86 416.66 431.86 417.1 426.51 417.1 426.51 418.1 296.825 418.1 296.825 418.355 273.39 418.355 273.39 418.35 151.735 418.35 151.735 418.355 136.64 418.355 136.64 418.1 5.35 418.1 5.35 417.1 0 417.1 0 416.66 8.81 416.66 8.81 412.6 0 412.6 0 412.16 5.35 412.16 5.35 411.16 136.64 411.16 136.64 410.92 296.825 410.92 296.825 411.16 426.51 411.16 426.51 412.16 431.86 412.16 ;
      RECT 410.37 0 411.815 5.88 ;
      RECT 386.37 0 386.81 5.88 ;
      POLYGON 431.86 475.6 0 475.6 0 475.16 5.35 475.16 5.35 474.16 126.6 474.16 126.6 474.205 130.02 474.205 130.02 474.16 136.64 474.16 136.64 473.92 293.995 473.92 293.995 474.205 297.415 474.205 297.415 474.16 426.51 474.16 426.51 475.16 431.86 475.16 ;
      POLYGON 244.225 484.88 242.97 484.88 242.97 481.56 237.41 481.56 237.41 484.88 236.845 484.88 236.845 481.16 244.225 481.16 ;
      RECT 310.07 0 311.195 5.88 ;
      POLYGON 431.86 106.13 426.51 106.13 426.51 108.855 419.095 108.855 419.095 108.85 280.11 108.85 280.11 111.175 139.41 111.175 139.41 108.85 119.9 108.85 119.9 108.855 5.35 108.855 5.35 106.13 0 106.13 0 103.975 147.285 103.975 147.285 108.405 147.325 108.405 147.325 108.815 221.88 108.815 221.88 108.82 278.505 108.82 278.505 103.975 431.86 103.975 ;
      POLYGON 287.455 484.88 285.23 484.88 285.23 481.56 279.67 481.56 279.67 484.88 276.59 484.88 276.59 481.16 287.455 481.16 ;
      RECT 277.57 0 278.51 5.88 ;
      POLYGON 431.86 277.6 423.05 277.6 423.05 281.66 431.86 281.66 431.86 282.1 426.51 282.1 426.51 283.1 296.825 283.1 296.825 283.355 273.39 283.355 273.39 283.35 151.735 283.35 151.735 283.355 136.64 283.355 136.64 283.1 5.35 283.1 5.35 282.1 0 282.1 0 281.66 8.81 281.66 8.81 277.6 0 277.6 0 277.16 5.35 277.16 5.35 276.16 136.64 276.16 136.64 275.92 296.825 275.92 296.825 276.16 426.51 276.16 426.51 277.16 431.86 277.16 ;
      POLYGON 176.795 484.88 175.4 484.88 175.4 481.56 169.84 481.56 169.84 484.88 167.185 484.88 167.185 481.56 161.625 481.56 161.625 484.88 158.83 484.88 158.83 481.16 176.795 481.16 ;
      POLYGON 195.86 5.88 185.435 5.88 185.435 0 189.86 0 189.86 4.94 195.42 4.94 195.42 0 195.86 0 ;
      POLYGON 431.86 28.55 277.69 28.55 277.69 27.745 254.33 27.745 254.33 32.68 207.265 32.68 207.265 30.605 173.39 30.605 173.39 28.045 147.01 28.045 147.01 28.55 0 28.55 0 28.425 118.155 28.425 118.155 28.43 136.35 28.43 136.35 25.595 121.53 25.595 121.53 25.59 15.335 25.59 15.335 25.585 8.84 25.585 8.84 22.855 119.265 22.855 119.265 23.375 289.265 23.375 289.265 23.385 312.425 23.385 312.425 22.855 423.02 22.855 423.02 25.585 416.525 25.585 416.525 25.59 308.73 25.59 308.73 25.595 289.265 25.595 289.265 28.43 312.425 28.43 312.425 28.425 431.86 28.425 ;
      RECT 241.445 0 242.55 5.88 ;
      POLYGON 33.725 484.88 32.09 484.88 32.09 481.56 26.53 481.56 26.53 484.88 25.965 484.88 25.965 481.16 33.725 481.16 ;
      POLYGON 431.86 403.6 423.05 403.6 423.05 407.66 431.86 407.66 431.86 408.1 426.51 408.1 426.51 409.1 296.825 409.1 296.825 409.355 273.39 409.355 273.39 409.35 151.735 409.35 151.735 409.355 136.64 409.355 136.64 409.1 5.35 409.1 5.35 408.1 0 408.1 0 407.66 8.81 407.66 8.81 403.6 0 403.6 0 403.16 5.35 403.16 5.35 402.16 136.64 402.16 136.64 401.92 296.825 401.92 296.825 402.16 426.51 402.16 426.51 403.16 431.86 403.16 ;
      POLYGON 431.86 268.6 423.05 268.6 423.05 272.66 431.86 272.66 431.86 273.1 426.51 273.1 426.51 274.1 296.825 274.1 296.825 274.355 273.39 274.355 273.39 274.35 151.735 274.35 151.735 274.355 136.64 274.355 136.64 274.1 5.35 274.1 5.35 273.1 0 273.1 0 272.66 8.81 272.66 8.81 268.6 0 268.6 0 268.16 5.35 268.16 5.35 267.16 136.64 267.16 136.64 266.92 296.825 266.92 296.825 267.16 426.51 267.16 426.51 268.16 431.86 268.16 ;
      POLYGON 426.51 34.63 424.215 34.63 424.215 34.62 308.845 34.62 308.845 34.625 308.73 34.625 308.73 34.64 277.69 34.64 277.69 31.275 312.425 31.275 312.425 31.27 416.525 31.27 416.525 31.275 426.51 31.275 ;
      POLYGON 431.86 259.6 423.05 259.6 423.05 263.66 431.86 263.66 431.86 264.1 426.51 264.1 426.51 265.1 296.825 265.1 296.825 265.355 273.39 265.355 273.39 265.35 151.735 265.35 151.735 265.355 136.64 265.355 136.64 265.1 5.35 265.1 5.35 264.1 0 264.1 0 263.66 8.81 263.66 8.81 259.6 0 259.6 0 259.16 5.35 259.16 5.35 258.16 136.64 258.16 136.64 257.92 296.825 257.92 296.825 258.16 426.51 258.16 426.51 259.16 431.86 259.16 ;
      POLYGON 431.86 385.6 423.05 385.6 423.05 389.66 431.86 389.66 431.86 390.1 426.51 390.1 426.51 391.1 296.825 391.1 296.825 391.355 273.39 391.355 273.39 391.35 151.735 391.35 151.735 391.355 136.64 391.355 136.64 391.1 5.35 391.1 5.35 390.1 0 390.1 0 389.66 8.81 389.66 8.81 385.6 0 385.6 0 385.16 5.35 385.16 5.35 384.16 136.64 384.16 136.64 383.92 296.825 383.92 296.825 384.16 426.51 384.16 426.51 385.16 431.86 385.16 ;
      POLYGON 117.135 484.88 116.57 484.88 116.57 481.56 111.01 481.56 111.01 484.88 108.545 484.88 108.545 481.16 117.135 481.16 ;
      POLYGON 431.86 40.48 308.845 40.48 308.845 40.485 308.73 40.485 308.73 40.49 289.265 40.49 289.265 47.86 311.67 47.86 311.67 47.855 362.45 47.855 362.45 47.85 362.73 47.85 362.73 47.855 416.45 47.855 416.45 47.85 426.51 47.85 426.51 47.855 431.86 47.855 431.86 50.6 422.69 50.6 422.69 50.585 308.845 50.585 308.845 50.595 308.745 50.595 308.745 50.6 286.195 50.6 286.195 53.42 211.025 53.42 211.025 57.735 308.845 57.735 308.845 57.745 431.86 57.745 431.86 59.9 425.275 59.9 425.275 59.895 292.035 59.895 292.035 58.205 207.86 58.205 207.86 49.58 173.425 49.58 173.425 53.5 147.11 53.5 147.11 58.94 133.58 58.94 133.58 59.95 121.53 59.95 121.53 59.9 0 59.9 0 57.745 15.335 57.745 15.335 57.735 119.955 57.735 119.955 57.745 139.42 57.745 139.42 50.6 121.53 50.6 121.53 50.59 10.965 50.59 10.965 50.595 10.865 50.595 10.865 50.6 0 50.6 0 47.855 5.35 47.855 5.35 47.85 10.85 47.85 10.85 47.855 119.955 47.855 119.955 47.86 143.925 47.86 143.925 38.54 173.39 38.54 173.39 33.44 147.405 33.44 147.405 35.14 140.61 35.14 140.61 40.49 121.53 40.49 121.53 40.485 15.335 40.485 15.335 40.48 0 40.48 0 38.26 15.335 38.26 15.335 38.255 117.845 38.255 117.845 38.26 139.42 38.26 139.42 34.63 121.53 34.63 121.53 34.62 10.965 34.62 10.965 34.625 10.85 34.625 10.85 34.63 5.35 34.63 5.35 31.275 15.335 31.275 15.335 31.27 118.155 31.27 118.155 31.275 147.01 31.275 147.01 33.145 174.02 33.145 174.02 39.22 147.285 39.22 147.285 43.19 207.265 43.19 207.265 37.24 254.33 37.24 254.33 45.545 209.005 45.545 209.005 52.38 257.43 52.38 257.43 47.79 277.69 47.79 277.69 44.93 288.96 44.93 288.96 38.26 314.015 38.26 314.015 38.255 416.525 38.255 416.525 38.26 431.86 38.26 ;
      POLYGON 431.86 376.6 423.05 376.6 423.05 380.66 431.86 380.66 431.86 381.1 426.51 381.1 426.51 382.1 296.825 382.1 296.825 382.355 273.39 382.355 273.39 382.35 151.735 382.35 151.735 382.355 136.64 382.355 136.64 382.1 5.35 382.1 5.35 381.1 0 381.1 0 380.66 8.81 380.66 8.81 376.6 0 376.6 0 376.16 5.35 376.16 5.35 375.16 136.64 375.16 136.64 374.92 296.825 374.92 296.825 375.16 426.51 375.16 426.51 376.16 431.86 376.16 ;
      POLYGON 345.285 484.88 343.29 484.88 343.29 481.56 337.73 481.56 337.73 484.88 337.165 484.88 337.165 481.16 345.285 481.16 ;
  END

END gf180mcu_fd_ip_sram__sram512x8m8wm1

END LIBRARY
