// //#############################################################################
// //# Function: Power isolation circuit                                         #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_isohi #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  iso,  // isolation signal
//     input  in,   // input
//     output out   // out = iso | in
// );
// 
//     assign out = iso | in;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
(* keep_hierarchy *)
module la_isohi (
    iso,
    in,
    out
);
  (* src = "generated" *)
  input in;
  wire in;
  (* src = "generated" *)
  input iso;
  wire iso;
  (* src = "generated" *)
  output out;
  wire out;
  gf180mcu_fd_sc_mcu9t5v0__or2_4 _0_ (
      .A1(in),
      .A2(iso),
      .Z (out)
  );
endmodule
