// //#############################################################################
// //# Function:  Reset synchronizer (async assert, sync deassert)               #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_rsync #(
//     parameter PROP = "DEFAULT"
// ) (
//     input clk,  // clock
//     input nrst_in,  // async reset input
//     output nrst_out  // async assert, sync deassert reset
// );
// 
//     localparam STAGES = 2;
//     localparam RND = 1;
// 
//     reg     [STAGES:0] sync_pipe;
//     integer            sync_delay;
// 
// `ifndef SYNTHESIS
//     always @(posedge clk) sync_delay <= {$random} % 2;
// `endif
// 
//     always @(posedge clk or negedge nrst_in)
//         if (!nrst_in) sync_pipe[STAGES:0] <= 'b0;
//         else sync_pipe[STAGES:0] <= {sync_pipe[STAGES-1:0], 1'b1};
// 
// `ifdef SYNTHESIS
//     assign nrst_out = sync_pipe[STAGES-1];
// `else
//     assign nrst_out = (|sync_delay & (|RND)) ? sync_pipe[STAGES] : sync_pipe[STAGES-1];
// `endif
// 
// endmodule

/* Generated by Yosys 0.38+92 (git sha1 84116c9a3, x86_64-conda-linux-gnu-cc 11.2.0 -fvisibility-inlines-hidden -fmessage-length=0 -march=nocona -mtune=haswell -ftree-vectorize -fPIC -fstack-protector-strong -fno-plt -O2 -ffunction-sections -fdebug-prefix-map=/root/conda-eda/conda-eda/workdir/conda-env/conda-bld/yosys_1708682838165/work=/usr/local/src/conda/yosys-0.38_93_g84116c9a3 -fdebug-prefix-map=/user/projekt_pia/miniconda3/envs/sc=/usr/local/src/conda-prefix -fPIC -Os -fno-merge-constants) */

module la_rsync(clk, nrst_in, nrst_out);
  wire _0_;
  input clk;
  wire clk;
  input nrst_in;
  wire nrst_in;
  output nrst_out;
  wire nrst_out;
  wire \sync_pipe[0] ;
  sky130_fd_sc_hdll__dfrtp_1 _1_ (
    .CLK(clk),
    .D(_0_),
    .Q(\sync_pipe[0] ),
    .RESET_B(nrst_in)
  );
  sky130_fd_sc_hdll__dfrtp_1 _2_ (
    .CLK(clk),
    .D(\sync_pipe[0] ),
    .Q(nrst_out),
    .RESET_B(nrst_in)
  );
  sky130_fd_sc_hdll__conb_1 _3_ (
    .HI(_0_)
  );
endmodule
