// //#############################################################################
// //# Function: Positive edge-triggered inverting static D-type flop-flop       #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_dffqn #(
//     parameter PROP = "DEFAULT"
// ) (
//     input d,
//     input clk,
//     output reg qn
// );
// 
//   always @(posedge clk) qn <= ~d;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_dffqn.v:10.1-20.10" *)
module la_dffqn (
    d,
    clk,
    qn
);
  (* src = "inputs/la_dffqn.v:18.3-18.34" *)
  wire _0_;
  wire _1_;
  (* src = "inputs/la_dffqn.v:14.11-14.14" *)
  input clk;
  wire clk;
  (* src = "inputs/la_dffqn.v:13.11-13.12" *)
  input d;
  wire d;
  (* src = "inputs/la_dffqn.v:15.16-15.18" *)
  output qn;
  wire qn;
  INVx2_ASAP7_75t_SL _2_ (
      .A(d),
      .Y(_0_)
  );
  INVx2_ASAP7_75t_SL _3_ (
      .A(_1_),
      .Y(qn)
  );
  (* src = "inputs/la_dffqn.v:18.3-18.34" *)
  DFFHQNx1_ASAP7_75t_SL _4_ (
      .CLK(clk),
      .D  (_0_),
      .QN (_1_)
  );
endmodule
