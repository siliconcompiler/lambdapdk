// //#############################################################################
// //# Function:  Positive edge-triggered static inverting D-type flop-flop with #
// //             async active low reset and scan input                          #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_sdffrqn #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      si,
//     input      se,
//     input      clk,
//     input      nreset,
//     output reg qn
// );
// 
//   always @(posedge clk or negedge nreset)
//     if (!nreset) qn <= 1'b1;
//     else qn <= se ? ~si : ~d;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_sdffrqn.v:11.1-26.10" *)
module la_sdffrqn (
    d,
    si,
    se,
    clk,
    nreset,
    qn
);
  (* src = "inputs/la_sdffrqn.v:22.3-24.30" *)
  wire _0_;
  wire _1_;
  (* src = "inputs/la_sdffrqn.v:17.16-17.19" *)
  input clk;
  wire clk;
  (* src = "inputs/la_sdffrqn.v:14.16-14.17" *)
  input d;
  wire d;
  (* src = "inputs/la_sdffrqn.v:18.16-18.22" *)
  input nreset;
  wire nreset;
  (* src = "inputs/la_sdffrqn.v:19.16-19.18" *)
  output qn;
  wire qn;
  (* src = "inputs/la_sdffrqn.v:16.16-16.18" *)
  input se;
  wire se;
  (* src = "inputs/la_sdffrqn.v:15.16-15.18" *)
  input si;
  wire si;
  gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2_ (
      .I0(d),
      .I1(si),
      .S (se),
      .Z (_1_)
  );
  gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3_ (
      .I (_1_),
      .ZN(_0_)
  );
  (* src = "inputs/la_sdffrqn.v:22.3-24.30" *)
  gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 _4_ (
      .CLK(clk),
      .D(_0_),
      .Q(qn),
      .SETN(nreset)
  );
endmodule
