// //#############################################################################
// //# Function: 2-Input Clock XOR Gate                                          #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_clkxor2 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a,
//     input  b,
//     output z
// );
// 
//     assign z = a ^ b;
// 
// endmodule

/* Generated by Yosys 0.40 (git sha1 a1bb0255d, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_clkxor2(a, b, z);
  input a;
  wire a;
  input b;
  wire b;
  output z;
  wire z;
  XOR2x1_ASAP7_75t_L _0_ (
    .A(b),
    .B(a),
    .Y(z)
  );
endmodule
