// //#############################################################################
// //# Function:  Positive edge-triggered static D-type flop-flop with async     #
// //#            active low reset.                                              #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_dffrq #(parameter PROP = "DEFAULT")   (
//     input      d,
//     input      clk,
//     input      nreset,
//     output reg q
//     );
// 
//    always @ (posedge clk or negedge nreset)
//      if(!nreset)
//        q <= 1'b0;
//      else
//        q <= d;
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_dffrq(d, clk, nreset, q);
  wire _0_;
  wire _1_;
  wire _2_;
  input clk;
  wire clk;
  input d;
  wire d;
  input nreset;
  wire nreset;
  output q;
  wire q;
  INVx2_ASAP7_75t_SL _3_ (
    .A(nreset),
    .Y(_1_)
  );
  INVx2_ASAP7_75t_SL _4_ (
    .A(_0_),
    .Y(q)
  );
  ASYNC_DFFHx1_ASAP7_75t_SL _5_ (
    .CLK(clk),
    .D(d),
    .QN(_0_),
    .RESET(_1_),
    .SET(_2_)
  );
  TIELOx1_ASAP7_75t_SL _6_ (
    .L(_2_)
  );
endmodule
