// //#############################################################################
// //# Function:  Positive edge-triggered static inverting D-type flop-flop with #
// //             async active low set.                                          #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_dffsqn #(parameter PROP = "DEFAULT")   (
//     input d,
//     input clk,
//     input nset,
//     output reg  qn
//     );
// 
//    always @ (posedge clk or negedge nset)
//      if(!nset)
//        qn <= 1'b0;
//      else
//        qn <= ~d;
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_dffsqn(d, clk, nset, qn);
  wire _0_;
  wire _1_;
  input clk;
  wire clk;
  input d;
  wire d;
  input nset;
  wire nset;
  output qn;
  wire qn;
  INV_X1 _2_ (
    .A(d),
    .ZN(_0_)
  );
  DFFR_X1 _3_ (
    .CK(clk),
    .D(_0_),
    .Q(qn),
    .QN(_1_),
    .RN(nset)
  );
endmodule
