// //#############################################################################
// //# Function:  Positive edge-triggered static D-type flop-flop with async     #
// //#            active low reset.                                              #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_dffrq #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      clk,
//     input      nreset,
//     output reg q
// );
// 
//     always @(posedge clk or negedge nreset)
//         if (!nreset) q <= 1'b0;
//         else q <= d;
// 
// endmodule

/* Generated by Yosys 0.40 (git sha1 a1bb0255d, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_dffrq(d, clk, nreset, q);
  wire _0_;
  wire _1_;
  input clk;
  wire clk;
  input d;
  wire d;
  input nreset;
  wire nreset;
  output q;
  wire q;
  INVx1_ASAP7_75t_R _2_ (
    .A(_0_),
    .Y(q)
  );
  DFFASRHQNx1_ASAP7_75t_R _3_ (
    .CLK(clk),
    .D(d),
    .QN(_0_),
    .RESETN(_1_),
    .SETN(nreset)
  );
  TIEHIx1_ASAP7_75t_R _4_ (
    .H(_1_)
  );
endmodule
