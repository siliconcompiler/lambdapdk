// //#############################################################################
// //# Function:  Positive edge-triggered static D-type flop-flop with async     #
// //#            active low preset.                                             #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_dffsq #(parameter PROP = "DEFAULT")   (
//     input      d,
//     input      clk,
//     input      nset,
//     output reg q
//     );
// 
//    always @ (posedge clk or negedge nset)
//      if(!nset)
//        q <= 1'b1;
//      else
//        q <= d;
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_dffsq(d, clk, nset, q);
  wire _0_;
  input clk;
  wire clk;
  input d;
  wire d;
  input nset;
  wire nset;
  output q;
  wire q;
  DFFS_X1 _1_ (
    .CK(clk),
    .D(d),
    .Q(q),
    .QN(_0_),
    .SN(nset)
  );
endmodule
