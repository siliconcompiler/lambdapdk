// //#############################################################################
// //# Function:  Positive edge-triggered static inverting D-type flop-flop with #
// //             async active low set.                                          #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_dffsqn #(parameter PROP = "DEFAULT")   (
//     input d,
//     input clk,
//     input nset,
//     output reg  qn
//     );
// 
//    always @ (posedge clk or negedge nset)
//      if(!nset)
//        qn <= 1'b0;
//      else
//        qn <= ~d;
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_dffsqn(d, clk, nset, qn);
  wire _0_;
  input clk;
  wire clk;
  input d;
  wire d;
  input nset;
  wire nset;
  output qn;
  wire qn;
  gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1_ (
    .I(d),
    .ZN(_0_)
  );
  gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 _2_ (
    .CLK(clk),
    .D(_0_),
    .Q(qn),
    .RN(nset)
  );
endmodule
