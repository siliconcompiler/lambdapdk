// //#############################################################################
// //# Function: Integrated "And" Clock Gating Cell (And)                        #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_clkicgand #(parameter PROP = "DEFAULT")  (
//    input  clk, // clock input
//    input  te, // test enable
//    input  en, // enable (from positive edge FF)
//    output eclk // enabled clock output
//    );
// 
//    reg 	  en_stable;
// 
//    always @ (clk or en or te)
//      if (~clk)
//        en_stable <= en | te;
// 
//    assign eclk =  clk & en_stable;
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_clkicgand(clk, te, en, eclk);
  wire _0_;
  input clk;
  wire clk;
  output eclk;
  wire eclk;
  input en;
  wire en;
  wire en_stable;
  input te;
  wire te;
  AND2_X1 _1_ (
    .A1(en_stable),
    .A2(clk),
    .ZN(eclk)
  );
  OR2_X2 _2_ (
    .A1(te),
    .A2(en),
    .ZN(_0_)
  );
  DLL_X1 _3_ (
    .D(_0_),
    .GN(clk),
    .Q(en_stable)
  );
endmodule
