// Source lambdapdk/gf180/libs/gf180mcu_fd_io/lef/5LM/gf180mcu_fd_io.lef

(* blackbox *)
module gf180mcu_fd_io__asig_5p0 (
    inout ASIG5V,
    inout DVDD,
    inout DVSS,
    inout VDD,
    inout VSS
);
endmodule

(* blackbox *)
module gf180mcu_fd_io__bi_24t (
    inout PAD,
    inout A,
    inout CS,
    inout IE,
    inout OE,
    inout PD,
    inout PU,
    inout SL,
    inout Y,
    inout DVDD,
    inout DVSS,
    inout VDD,
    inout VSS
);
endmodule

(* blackbox *)
module gf180mcu_fd_io__bi_t (
    inout PAD,
    inout A,
    inout CS,
    inout IE,
    inout OE,
    inout PD,
    inout PDRV0,
    inout PDRV1,
    inout PU,
    inout SL,
    inout Y,
    inout DVDD,
    inout DVSS,
    inout VDD,
    inout VSS
);
endmodule

(* blackbox *)
module gf180mcu_fd_io__brk2 (
    inout VSS
);
endmodule

(* blackbox *)
module gf180mcu_fd_io__brk5 (
    inout VSS
);
endmodule

(* blackbox *)
module gf180mcu_fd_io__cor (
    inout DVDD,
    inout DVSS,
    inout VDD,
    inout VSS
);
endmodule

(* blackbox *)
module gf180mcu_fd_io__dvdd (
    inout DVDD,
    inout DVSS,
    inout VSS
);
endmodule

(* blackbox *)
module gf180mcu_fd_io__dvss (
    inout DVSS,
    inout DVDD,
    inout VDD
);
endmodule

(* blackbox *)
module gf180mcu_fd_io__fill1 (
    inout DVDD,
    inout DVSS,
    inout VDD,
    inout VSS
);
endmodule

(* blackbox *)
module gf180mcu_fd_io__fill5 (
    inout DVDD,
    inout DVSS,
    inout VDD,
    inout VSS
);
endmodule

(* blackbox *)
module gf180mcu_fd_io__fill10 (
    inout DVDD,
    inout DVSS,
    inout VDD,
    inout VSS
);
endmodule

(* blackbox *)
module gf180mcu_fd_io__fillnc (
    inout DVDD,
    inout DVSS,
    inout VDD,
    inout VSS
);
endmodule

(* blackbox *)
module gf180mcu_fd_io__in_c (
    inout PAD,
    inout PD,
    inout PU,
    inout Y,
    inout DVDD,
    inout DVSS,
    inout VDD,
    inout VSS
);
endmodule

(* blackbox *)
module gf180mcu_fd_io__in_s (
    inout PAD,
    inout PD,
    inout PU,
    inout Y,
    inout DVDD,
    inout DVSS,
    inout VDD,
    inout VSS
);
endmodule
