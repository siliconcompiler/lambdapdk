// //#############################################################################
// //# Function: 3-Input one-hot mux                                             #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_dmux3
//   #(parameter PROP = "DEFAULT")
//    (
//     input  sel0,
//     input  sel1,
//     input  sel2,
//     input  in0,
//     input  in1,
//     input  in2,
//     output out
//     );
// 
//    assign out = (sel0 & in0) |
// 		(sel1 & in1) |
// 		(sel2 & in2);
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_dmux3(sel0, sel1, sel2, in0, in1, in2, out);
  wire _0_;
  input in0;
  wire in0;
  input in1;
  wire in1;
  input in2;
  wire in2;
  output out;
  wire out;
  input sel0;
  wire sel0;
  input sel1;
  wire sel1;
  input sel2;
  wire sel2;
  sky130_fd_sc_hd__a222oi_1 _1_ (
    .A1(in0),
    .A2(sel0),
    .B1(in1),
    .B2(sel1),
    .C1(in2),
    .C2(sel2),
    .Y(_0_)
  );
  sky130_fd_sc_hd__inv_1 _2_ (
    .A(_0_),
    .Y(out)
  );
endmodule
