VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO fakepll7
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 100 BY 100 ;
  SYMMETRY X Y ;

  #-----------------------------------------------------------------------------
  # Power Pins (Layer M5) - Vertical Stripes
  # Spanning y=0 to y=100
  #-----------------------------------------------------------------------------
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
      RECT 20.000 0.000 21.000 100.000 ; 
      RECT 25.000 0.000 26.000 100.000 ; 
    END
  END VDDA

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
      RECT 40.000 0.000 41.000 100.000 ;
      RECT 45.000 0.000 46.000 100.000 ;
    END
  END VDD

  PIN VDD2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
      RECT 60.000 0.000 61.000 100.000 ;
      RECT 65.000 0.000 66.000 100.000 ;
    END
  END VDD2

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
      RECT 80.000 0.000 81.000 100.000 ;
      RECT 85.000 0.000 86.000 100.000 ;
    END
  END VSS

  #-----------------------------------------------------------------------------
  # INPUT PINS (Left Side) - Layer M4
  # x coordinates: 0.000 to 1.000
  #-----------------------------------------------------------------------------

  # --- Reference Clocks ---
  PIN clkin[0]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 1.000 1.000 1.024 ; END
  END clkin[0]
  PIN clkin[1]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 1.450 1.000 1.474 ; END
  END clkin[1]

  # --- Feedback Input ---
  PIN clkfbin
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 1.900 1.000 1.924 ; END
  END clkfbin

  # --- Standard Controls ---
  PIN reset
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 2.350 1.000 2.374 ; END
  END reset
  PIN en
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 2.800 1.000 2.824 ; END
  END en
  PIN bypass
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 3.250 1.000 3.274 ; END
  END bypass
  PIN clksel[0]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 3.700 1.000 3.724 ; END
  END clksel[0]

  # --- Clock Enables (8 bits) ---
  PIN clken[0]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 4.150 1.000 4.174 ; END
  END clken[0]
  PIN clken[1]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 4.600 1.000 4.624 ; END
  END clken[1]
  PIN clken[2]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 5.050 1.000 5.074 ; END
  END clken[2]
  PIN clken[3]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 5.500 1.000 5.524 ; END
  END clken[3]
  PIN clken[4]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 5.950 1.000 5.974 ; END
  END clken[4]
  PIN clken[5]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 6.400 1.000 6.424 ; END
  END clken[5]
  PIN clken[6]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 6.850 1.000 6.874 ; END
  END clken[6]
  PIN clken[7]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 7.300 1.000 7.324 ; END
  END clken[7]

  # --- Input Divider (8 bits) ---
  PIN divin[0]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 7.750 1.000 7.774 ; END
  END divin[0]
  PIN divin[1]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 8.200 1.000 8.224 ; END
  END divin[1]
  PIN divin[2]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 8.650 1.000 8.674 ; END
  END divin[2]
  PIN divin[3]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 9.100 1.000 9.124 ; END
  END divin[3]
  PIN divin[4]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 9.550 1.000 9.574 ; END
  END divin[4]
  PIN divin[5]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 10.000 1.000 10.024 ; END
  END divin[5]
  PIN divin[6]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 10.450 1.000 10.474 ; END
  END divin[6]
  PIN divin[7]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 10.900 1.000 10.924 ; END
  END divin[7]

  # --- Feedback Divider (16 bits) ---
  PIN divfb[0]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 11.350 1.000 11.374 ; END
  END divfb[0]
  PIN divfb[1]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 11.800 1.000 11.824 ; END
  END divfb[1]
  PIN divfb[2]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 12.250 1.000 12.274 ; END
  END divfb[2]
  PIN divfb[3]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 12.700 1.000 12.724 ; END
  END divfb[3]
  PIN divfb[4]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 13.150 1.000 13.174 ; END
  END divfb[4]
  PIN divfb[5]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 13.600 1.000 13.624 ; END
  END divfb[5]
  PIN divfb[6]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 14.050 1.000 14.074 ; END
  END divfb[6]
  PIN divfb[7]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 14.500 1.000 14.524 ; END
  END divfb[7]
  PIN divfb[8]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 14.950 1.000 14.974 ; END
  END divfb[8]
  PIN divfb[9]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 15.400 1.000 15.424 ; END
  END divfb[9]
  PIN divfb[10]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 15.850 1.000 15.874 ; END
  END divfb[10]
  PIN divfb[11]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 16.300 1.000 16.324 ; END
  END divfb[11]
  PIN divfb[12]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 16.750 1.000 16.774 ; END
  END divfb[12]
  PIN divfb[13]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 17.200 1.000 17.224 ; END
  END divfb[13]
  PIN divfb[14]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 17.650 1.000 17.674 ; END
  END divfb[14]
  PIN divfb[15]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 18.100 1.000 18.124 ; END
  END divfb[15]

  # --- Fractional Divider (8 bits) ---
  PIN divfrac[0]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 18.550 1.000 18.574 ; END
  END divfrac[0]
  PIN divfrac[1]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 19.000 1.000 19.024 ; END
  END divfrac[1]
  PIN divfrac[2]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 19.450 1.000 19.474 ; END
  END divfrac[2]
  PIN divfrac[3]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 19.900 1.000 19.924 ; END
  END divfrac[3]
  PIN divfrac[4]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 20.350 1.000 20.374 ; END
  END divfrac[4]
  PIN divfrac[5]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 20.800 1.000 20.824 ; END
  END divfrac[5]
  PIN divfrac[6]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 21.250 1.000 21.274 ; END
  END divfrac[6]
  PIN divfrac[7]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 21.700 1.000 21.724 ; END
  END divfrac[7]

  # --- Output Dividers (64 bits) ---
  PIN divout[0]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 22.150 1.000 22.174 ; END
  END divout[0]
  PIN divout[1]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 22.600 1.000 22.624 ; END
  END divout[1]
  PIN divout[2]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 23.050 1.000 23.074 ; END
  END divout[2]
  PIN divout[3]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 23.500 1.000 23.524 ; END
  END divout[3]
  PIN divout[4]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 23.950 1.000 23.974 ; END
  END divout[4]
  PIN divout[5]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 24.400 1.000 24.424 ; END
  END divout[5]
  PIN divout[6]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 24.850 1.000 24.874 ; END
  END divout[6]
  PIN divout[7]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 25.300 1.000 25.324 ; END
  END divout[7]
  PIN divout[8]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 25.750 1.000 25.774 ; END
  END divout[8]
  PIN divout[9]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 26.200 1.000 26.224 ; END
  END divout[9]
  PIN divout[10]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 26.650 1.000 26.674 ; END
  END divout[10]
  PIN divout[11]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 27.100 1.000 27.124 ; END
  END divout[11]
  PIN divout[12]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 27.550 1.000 27.574 ; END
  END divout[12]
  PIN divout[13]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 28.000 1.000 28.024 ; END
  END divout[13]
  PIN divout[14]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 28.450 1.000 28.474 ; END
  END divout[14]
  PIN divout[15]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 28.900 1.000 28.924 ; END
  END divout[15]
  PIN divout[16]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 29.350 1.000 29.374 ; END
  END divout[16]
  PIN divout[17]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 29.800 1.000 29.824 ; END
  END divout[17]
  PIN divout[18]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 30.250 1.000 30.274 ; END
  END divout[18]
  PIN divout[19]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 30.700 1.000 30.724 ; END
  END divout[19]
  PIN divout[20]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 31.150 1.000 31.174 ; END
  END divout[20]
  PIN divout[21]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 31.600 1.000 31.624 ; END
  END divout[21]
  PIN divout[22]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 32.050 1.000 32.074 ; END
  END divout[22]
  PIN divout[23]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 32.500 1.000 32.524 ; END
  END divout[23]
  PIN divout[24]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 32.950 1.000 32.974 ; END
  END divout[24]
  PIN divout[25]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 33.400 1.000 33.424 ; END
  END divout[25]
  PIN divout[26]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 33.850 1.000 33.874 ; END
  END divout[26]
  PIN divout[27]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 34.300 1.000 34.324 ; END
  END divout[27]
  PIN divout[28]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 34.750 1.000 34.774 ; END
  END divout[28]
  PIN divout[29]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 35.200 1.000 35.224 ; END
  END divout[29]
  PIN divout[30]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 35.650 1.000 35.674 ; END
  END divout[30]
  PIN divout[31]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 36.100 1.000 36.124 ; END
  END divout[31]
  PIN divout[32]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 36.550 1.000 36.574 ; END
  END divout[32]
  PIN divout[33]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 37.000 1.000 37.024 ; END
  END divout[33]
  PIN divout[34]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 37.450 1.000 37.474 ; END
  END divout[34]
  PIN divout[35]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 37.900 1.000 37.924 ; END
  END divout[35]
  PIN divout[36]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 38.350 1.000 38.374 ; END
  END divout[36]
  PIN divout[37]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 38.800 1.000 38.824 ; END
  END divout[37]
  PIN divout[38]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 39.250 1.000 39.274 ; END
  END divout[38]
  PIN divout[39]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 39.700 1.000 39.724 ; END
  END divout[39]
  PIN divout[40]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 40.150 1.000 40.174 ; END
  END divout[40]
  PIN divout[41]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 40.600 1.000 40.624 ; END
  END divout[41]
  PIN divout[42]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 41.050 1.000 41.074 ; END
  END divout[42]
  PIN divout[43]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 41.500 1.000 41.524 ; END
  END divout[43]
  PIN divout[44]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 41.950 1.000 41.974 ; END
  END divout[44]
  PIN divout[45]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 42.400 1.000 42.424 ; END
  END divout[45]
  PIN divout[46]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 42.850 1.000 42.874 ; END
  END divout[46]
  PIN divout[47]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 43.300 1.000 43.324 ; END
  END divout[47]
  PIN divout[48]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 43.750 1.000 43.774 ; END
  END divout[48]
  PIN divout[49]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 44.200 1.000 44.224 ; END
  END divout[49]
  PIN divout[50]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 44.650 1.000 44.674 ; END
  END divout[50]
  PIN divout[51]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 45.100 1.000 45.124 ; END
  END divout[51]
  PIN divout[52]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 45.550 1.000 45.574 ; END
  END divout[52]
  PIN divout[53]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 46.000 1.000 46.024 ; END
  END divout[53]
  PIN divout[54]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 46.450 1.000 46.474 ; END
  END divout[54]
  PIN divout[55]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 46.900 1.000 46.924 ; END
  END divout[55]
  PIN divout[56]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 47.350 1.000 47.374 ; END
  END divout[56]
  PIN divout[57]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 47.800 1.000 47.824 ; END
  END divout[57]
  PIN divout[58]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 48.250 1.000 48.274 ; END
  END divout[58]
  PIN divout[59]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 48.700 1.000 48.724 ; END
  END divout[59]
  PIN divout[60]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 49.150 1.000 49.174 ; END
  END divout[60]
  PIN divout[61]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 49.600 1.000 49.624 ; END
  END divout[61]
  PIN divout[62]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 50.050 1.000 50.074 ; END
  END divout[62]
  PIN divout[63]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 50.500 1.000 50.524 ; END
  END divout[63]

  # --- Phase Shift (64 bits) ---
  PIN phase[0]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 50.950 1.000 50.974 ; END
  END phase[0]
  PIN phase[1]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 51.400 1.000 51.424 ; END
  END phase[1]
  PIN phase[2]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 51.850 1.000 51.874 ; END
  END phase[2]
  PIN phase[3]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 52.300 1.000 52.324 ; END
  END phase[3]
  PIN phase[4]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 52.750 1.000 52.774 ; END
  END phase[4]
  PIN phase[5]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 53.200 1.000 53.224 ; END
  END phase[5]
  PIN phase[6]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 53.650 1.000 53.674 ; END
  END phase[6]
  PIN phase[7]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 54.100 1.000 54.124 ; END
  END phase[7]
  PIN phase[8]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 54.550 1.000 54.574 ; END
  END phase[8]
  PIN phase[9]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 55.000 1.000 55.024 ; END
  END phase[9]
  PIN phase[10]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 55.450 1.000 55.474 ; END
  END phase[10]
  PIN phase[11]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 55.900 1.000 55.924 ; END
  END phase[11]
  PIN phase[12]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 56.350 1.000 56.374 ; END
  END phase[12]
  PIN phase[13]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 56.800 1.000 56.824 ; END
  END phase[13]
  PIN phase[14]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 57.250 1.000 57.274 ; END
  END phase[14]
  PIN phase[15]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 57.700 1.000 57.724 ; END
  END phase[15]
  PIN phase[16]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 58.150 1.000 58.174 ; END
  END phase[16]
  PIN phase[17]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 58.600 1.000 58.624 ; END
  END phase[17]
  PIN phase[18]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 59.050 1.000 59.074 ; END
  END phase[18]
  PIN phase[19]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 59.500 1.000 59.524 ; END
  END phase[19]
  PIN phase[20]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 59.950 1.000 59.974 ; END
  END phase[20]
  PIN phase[21]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 60.400 1.000 60.424 ; END
  END phase[21]
  PIN phase[22]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 60.850 1.000 60.874 ; END
  END phase[22]
  PIN phase[23]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 61.300 1.000 61.324 ; END
  END phase[23]
  PIN phase[24]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 61.750 1.000 61.774 ; END
  END phase[24]
  PIN phase[25]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 62.200 1.000 62.224 ; END
  END phase[25]
  PIN phase[26]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 62.650 1.000 62.674 ; END
  END phase[26]
  PIN phase[27]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 63.100 1.000 63.124 ; END
  END phase[27]
  PIN phase[28]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 63.550 1.000 63.574 ; END
  END phase[28]
  PIN phase[29]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 64.000 1.000 64.024 ; END
  END phase[29]
  PIN phase[30]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 64.450 1.000 64.474 ; END
  END phase[30]
  PIN phase[31]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 64.900 1.000 64.924 ; END
  END phase[31]
  PIN phase[32]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 65.350 1.000 65.374 ; END
  END phase[32]
  PIN phase[33]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 65.800 1.000 65.824 ; END
  END phase[33]
  PIN phase[34]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 66.250 1.000 66.274 ; END
  END phase[34]
  PIN phase[35]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 66.700 1.000 66.724 ; END
  END phase[35]
  PIN phase[36]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 67.150 1.000 67.174 ; END
  END phase[36]
  PIN phase[37]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 67.600 1.000 67.624 ; END
  END phase[37]
  PIN phase[38]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 68.050 1.000 68.074 ; END
  END phase[38]
  PIN phase[39]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 68.500 1.000 68.524 ; END
  END phase[39]
  PIN phase[40]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 68.950 1.000 68.974 ; END
  END phase[40]
  PIN phase[41]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 69.400 1.000 69.424 ; END
  END phase[41]
  PIN phase[42]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 69.850 1.000 69.874 ; END
  END phase[42]
  PIN phase[43]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 70.300 1.000 70.324 ; END
  END phase[43]
  PIN phase[44]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 70.750 1.000 70.774 ; END
  END phase[44]
  PIN phase[45]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 71.200 1.000 71.224 ; END
  END phase[45]
  PIN phase[46]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 71.650 1.000 71.674 ; END
  END phase[46]
  PIN phase[47]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 72.100 1.000 72.124 ; END
  END phase[47]
  PIN phase[48]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 72.550 1.000 72.574 ; END
  END phase[48]
  PIN phase[49]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 73.000 1.000 73.024 ; END
  END phase[49]
  PIN phase[50]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 73.450 1.000 73.474 ; END
  END phase[50]
  PIN phase[51]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 73.900 1.000 73.924 ; END
  END phase[51]
  PIN phase[52]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 74.350 1.000 74.374 ; END
  END phase[52]
  PIN phase[53]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 74.800 1.000 74.824 ; END
  END phase[53]
  PIN phase[54]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 75.250 1.000 75.274 ; END
  END phase[54]
  PIN phase[55]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 75.700 1.000 75.724 ; END
  END phase[55]
  PIN phase[56]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 76.150 1.000 76.174 ; END
  END phase[56]
  PIN phase[57]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 76.600 1.000 76.624 ; END
  END phase[57]
  PIN phase[58]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 77.050 1.000 77.074 ; END
  END phase[58]
  PIN phase[59]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 77.500 1.000 77.524 ; END
  END phase[59]
  PIN phase[60]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 77.950 1.000 77.974 ; END
  END phase[60]
  PIN phase[61]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 78.400 1.000 78.424 ; END
  END phase[61]
  PIN phase[62]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 78.850 1.000 78.874 ; END
  END phase[62]
  PIN phase[63]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 79.300 1.000 79.324 ; END
  END phase[63]

  # --- Controls (32 bits) ---
  PIN ctrl[0]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 79.750 1.000 79.774 ; END
  END ctrl[0]
  PIN ctrl[1]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 80.200 1.000 80.224 ; END
  END ctrl[1]
  PIN ctrl[2]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 80.650 1.000 80.674 ; END
  END ctrl[2]
  PIN ctrl[3]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 81.100 1.000 81.124 ; END
  END ctrl[3]
  PIN ctrl[4]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 81.550 1.000 81.574 ; END
  END ctrl[4]
  PIN ctrl[5]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 82.000 1.000 82.024 ; END
  END ctrl[5]
  PIN ctrl[6]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 82.450 1.000 82.474 ; END
  END ctrl[6]
  PIN ctrl[7]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 82.900 1.000 82.924 ; END
  END ctrl[7]
  PIN ctrl[8]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 83.350 1.000 83.374 ; END
  END ctrl[8]
  PIN ctrl[9]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 83.800 1.000 83.824 ; END
  END ctrl[9]
  PIN ctrl[10]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 84.250 1.000 84.274 ; END
  END ctrl[10]
  PIN ctrl[11]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 84.700 1.000 84.724 ; END
  END ctrl[11]
  PIN ctrl[12]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 85.150 1.000 85.174 ; END
  END ctrl[12]
  PIN ctrl[13]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 85.600 1.000 85.624 ; END
  END ctrl[13]
  PIN ctrl[14]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 86.050 1.000 86.074 ; END
  END ctrl[14]
  PIN ctrl[15]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 86.500 1.000 86.524 ; END
  END ctrl[15]
  PIN ctrl[16]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 86.950 1.000 86.974 ; END
  END ctrl[16]
  PIN ctrl[17]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 87.400 1.000 87.424 ; END
  END ctrl[17]
  PIN ctrl[18]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 87.850 1.000 87.874 ; END
  END ctrl[18]
  PIN ctrl[19]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 88.300 1.000 88.324 ; END
  END ctrl[19]
  PIN ctrl[20]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 88.750 1.000 88.774 ; END
  END ctrl[20]
  PIN ctrl[21]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 89.200 1.000 89.224 ; END
  END ctrl[21]
  PIN ctrl[22]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 89.650 1.000 89.674 ; END
  END ctrl[22]
  PIN ctrl[23]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 90.100 1.000 90.124 ; END
  END ctrl[23]
  PIN ctrl[24]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 90.550 1.000 90.574 ; END
  END ctrl[24]
  PIN ctrl[25]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 91.000 1.000 91.024 ; END
  END ctrl[25]
  PIN ctrl[26]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 91.450 1.000 91.474 ; END
  END ctrl[26]
  PIN ctrl[27]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 91.900 1.000 91.924 ; END
  END ctrl[27]
  PIN ctrl[28]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 92.350 1.000 92.374 ; END
  END ctrl[28]
  PIN ctrl[29]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 92.800 1.000 92.824 ; END
  END ctrl[29]
  PIN ctrl[30]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 93.250 1.000 93.274 ; END
  END ctrl[30]
  PIN ctrl[31]
    DIRECTION INPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 0.000 93.700 1.000 93.724 ; END
  END ctrl[31]

  #-----------------------------------------------------------------------------
  # OUTPUT PINS (Right Side) - Layer M4
  # x coordinates: 99.000 to 100.000
  #-----------------------------------------------------------------------------

  # --- Output Clocks (8 bits) ---
  PIN clkout[0]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 1.000 100.000 1.024 ; END
  END clkout[0]
  PIN clkout[1]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 3.000 100.000 3.024 ; END
  END clkout[1]
  PIN clkout[2]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 5.000 100.000 5.024 ; END
  END clkout[2]
  PIN clkout[3]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 7.000 100.000 7.024 ; END
  END clkout[3]
  PIN clkout[4]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 9.000 100.000 9.024 ; END
  END clkout[4]
  PIN clkout[5]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 11.000 100.000 11.024 ; END
  END clkout[5]
  PIN clkout[6]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 13.000 100.000 13.024 ; END
  END clkout[6]
  PIN clkout[7]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 15.000 100.000 15.024 ; END
  END clkout[7]

  # --- Feedback/VCO ---
  PIN clkfbout
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 17.000 100.000 17.024 ; END
  END clkfbout
  PIN clkvco
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 19.000 100.000 19.024 ; END
  END clkvco

  # --- Locks ---
  PIN freqlock
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 21.000 100.000 21.024 ; END
  END freqlock
  PIN phaselock
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 23.000 100.000 23.024 ; END
  END phaselock

  # --- Status (32 bits) ---
  PIN status[0]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 25.000 100.000 25.024 ; END
  END status[0]
  PIN status[1]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 27.000 100.000 27.024 ; END
  END status[1]
  PIN status[2]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 29.000 100.000 29.024 ; END
  END status[2]
  PIN status[3]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 31.000 100.000 31.024 ; END
  END status[3]
  PIN status[4]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 33.000 100.000 33.024 ; END
  END status[4]
  PIN status[5]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 35.000 100.000 35.024 ; END
  END status[5]
  PIN status[6]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 37.000 100.000 37.024 ; END
  END status[6]
  PIN status[7]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 39.000 100.000 39.024 ; END
  END status[7]
  PIN status[8]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 41.000 100.000 41.024 ; END
  END status[8]
  PIN status[9]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 43.000 100.000 43.024 ; END
  END status[9]
  PIN status[10]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 45.000 100.000 45.024 ; END
  END status[10]
  PIN status[11]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 47.000 100.000 47.024 ; END
  END status[11]
  PIN status[12]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 49.000 100.000 49.024 ; END
  END status[12]
  PIN status[13]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 51.000 100.000 51.024 ; END
  END status[13]
  PIN status[14]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 53.000 100.000 53.024 ; END
  END status[14]
  PIN status[15]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 55.000 100.000 55.024 ; END
  END status[15]
  PIN status[16]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 57.000 100.000 57.024 ; END
  END status[16]
  PIN status[17]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 59.000 100.000 59.024 ; END
  END status[17]
  PIN status[18]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 61.000 100.000 61.024 ; END
  END status[18]
  PIN status[19]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 63.000 100.000 63.024 ; END
  END status[19]
  PIN status[20]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 65.000 100.000 65.024 ; END
  END status[20]
  PIN status[21]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 67.000 100.000 67.024 ; END
  END status[21]
  PIN status[22]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 69.000 100.000 69.024 ; END
  END status[22]
  PIN status[23]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 71.000 100.000 71.024 ; END
  END status[23]
  PIN status[24]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 73.000 100.000 73.024 ; END
  END status[24]
  PIN status[25]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 75.000 100.000 75.024 ; END
  END status[25]
  PIN status[26]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 77.000 100.000 77.024 ; END
  END status[26]
  PIN status[27]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 79.000 100.000 79.024 ; END
  END status[27]
  PIN status[28]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 81.000 100.000 81.024 ; END
  END status[28]
  PIN status[29]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 83.000 100.000 83.024 ; END
  END status[29]
  PIN status[30]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 85.000 100.000 85.024 ; END
  END status[30]
  PIN status[31]
    DIRECTION OUTPUT ; USE SIGNAL ; PORT LAYER M4 ; RECT 99.000 87.000 100.000 87.024 ; END
  END status[31]

END fakepll7
