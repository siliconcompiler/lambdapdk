// //#############################################################################
// //# Function: Positive edge-triggered static D-type flop-flop with scan input #
// //#                                                                           #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_sdffq #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      si,
//     input      se,
//     input      clk,
//     output reg q
// );
// 
//     always @(posedge clk) q <= se ? si : d;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
module la_sdffq (
    d,
    si,
    se,
    clk,
    q
);
  (* src = "generated" *)
  wire _0_;
  wire _1_;
  wire _2_;
  wire _3_;
  (* src = "generated" *)
  input clk;
  wire clk;
  (* src = "generated" *)
  input d;
  wire d;
  (* src = "generated" *)
  output q;
  wire q;
  (* src = "generated" *)
  input se;
  wire se;
  (* src = "generated" *)
  input si;
  wire si;
  INVx1_ASAP7_75t_L _4_ (
      .A(se),
      .Y(_2_)
  );
  AND2x2_ASAP7_75t_L _5_ (
      .A(si),
      .B(se),
      .Y(_3_)
  );
  AO21x1_ASAP7_75t_L _6_ (
      .A1(d),
      .A2(_2_),
      .B (_3_),
      .Y (_0_)
  );
  INVx1_ASAP7_75t_L _7_ (
      .A(_1_),
      .Y(q)
  );
  (* src = "generated" *)
  DFFHQNx1_ASAP7_75t_L _8_ (
      .CLK(clk),
      .D  (_0_),
      .QN (_1_)
  );
endmodule
