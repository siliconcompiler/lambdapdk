// //#############################################################################
// //# Function: Dual data rate input buffer                                     #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_iddr #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      clk,      // clock
//     input      in,       // data input sampled on both edges of clock
//     output reg outrise,  // rising edge sample
//     output reg outfall   // falling edge sample
// );
// 
//     // Negedge Sample
//     always @(negedge clk) outfall <= in;
// 
//     // Posedge Sample
//     reg inrise;
//     always @(posedge clk) inrise <= in;
// 
//     // Posedge Latch (for hold)
//     always @(clk or inrise) if (~clk) outrise <= inrise;
// 
// endmodule

/* Generated by Yosys 0.41 (git sha1 c1ad37779, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_iddr(clk, in, outrise, outfall);
  wire _0_;
  input clk;
  wire clk;
  input in;
  wire in;
  wire inrise;
  output outfall;
  wire outfall;
  output outrise;
  wire outrise;
  gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1_ (
    .I(clk),
    .ZN(_0_)
  );
  gf180mcu_fd_sc_mcu9t5v0__latq_1 _2_ (
    .D(inrise),
    .E(_0_),
    .Q(outrise)
  );
  gf180mcu_fd_sc_mcu9t5v0__dffq_2 _3_ (
    .CLK(clk),
    .D(in),
    .Q(inrise)
  );
  gf180mcu_fd_sc_mcu9t5v0__dffnq_2 _4_ (
    .CLKN(clk),
    .D(in),
    .Q(outfall)
  );
endmodule
