// //#############################################################################
// //# Function: And-Or (ao221) Gate                                             #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_ao221 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  a0,
//     input  a1,
//     input  b0,
//     input  b1,
//     input  c0,
//     output z
// );
// 
//     assign z = (a0 & a1) | (b0 & b1) | (c0);
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
(* keep_hierarchy *)
module la_ao221 (
    a0,
    a1,
    b0,
    b1,
    c0,
    z
);
  wire _0_;
  (* src = "generated" *)
  input a0;
  wire a0;
  (* src = "generated" *)
  input a1;
  wire a1;
  (* src = "generated" *)
  input b0;
  wire b0;
  (* src = "generated" *)
  input b1;
  wire b1;
  (* src = "generated" *)
  input c0;
  wire c0;
  (* src = "generated" *)
  output z;
  wire z;
  gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _1_ (
      .A1(a1),
      .A2(a0),
      .B1(b1),
      .B2(b0),
      .C (c0),
      .ZN(_0_)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_2 _2_ (
      .I (_0_),
      .ZN(z)
  );
endmodule
