// Source ../.sc/cache/ihp130-62c1d640dc1c91f5-1d3cde26ed72789c/ihp-sg13g2/libs.ref/sg13g2_io/lef/sg13g2_io.lef

(* blackbox *)
module sg13g2_Corner (
    inout iovdd,
    inout iovss,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_Filler200 (
    inout iovdd,
    inout iovss,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_Filler400 (
    inout iovdd,
    inout iovss,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_Filler1000 (
    inout iovdd,
    inout iovss,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_Filler2000 (
    inout iovdd,
    inout iovss,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_Filler4000 (
    inout iovdd,
    inout iovss,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_Filler10000 (
    inout iovdd,
    inout iovss,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadIn (
    inout iovdd,
    inout iovss,
    output p2c,
    inout pad,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadOut4mA (
    input c2p,
    inout iovdd,
    inout iovss,
    inout pad,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadOut16mA (
    input c2p,
    inout iovdd,
    inout iovss,
    inout pad,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadOut30mA (
    input c2p,
    inout iovdd,
    inout iovss,
    inout pad,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadTriOut4mA (
    input c2p,
    input c2p_en,
    inout iovdd,
    inout iovss,
    inout pad,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadTriOut16mA (
    input c2p,
    input c2p_en,
    inout iovdd,
    inout iovss,
    inout pad,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadTriOut30mA (
    input c2p,
    input c2p_en,
    inout iovdd,
    inout iovss,
    inout pad,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadInOut4mA (
    input c2p,
    input c2p_en,
    inout iovdd,
    inout iovss,
    output p2c,
    inout pad,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadInOut16mA (
    input c2p,
    input c2p_en,
    inout iovdd,
    inout iovss,
    output p2c,
    inout pad,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadInOut30mA (
    input c2p,
    input c2p_en,
    inout iovdd,
    inout iovss,
    output p2c,
    inout pad,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadAnalog (
    inout iovdd,
    inout iovss,
    inout pad,
    inout padres,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadIOVss (
    inout iovdd,
    inout iovss,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadIOVdd (
    inout iovdd,
    inout iovss,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadVss (
    inout iovdd,
    inout iovss,
    inout vdd,
    inout vss
);
endmodule

(* blackbox *)
module sg13g2_IOPadVdd (
    inout iovdd,
    inout iovss,
    inout vdd,
    inout vss
);
endmodule
