// //#############################################################################
// //# Function:  Positive edge-triggered static inverting D-type flop-flop with #
// //             async active low reset.                                        #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_dffrqn #(parameter PROP = "DEFAULT")   (
//     input      d,
//     input      clk,
//     input      nreset,
//     output reg qn
//     );
// 
//    always @ (posedge clk or negedge nreset)
//      if(!nreset)
//        qn <= 1'b1;
//      else
//        qn <= ~d;
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_dffrqn(d, clk, nreset, qn);
  wire _0_;
  input clk;
  wire clk;
  input d;
  wire d;
  input nreset;
  wire nreset;
  output qn;
  wire qn;
  gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1_ (
    .I(d),
    .ZN(_0_)
  );
  gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 _2_ (
    .CLK(clk),
    .D(_0_),
    .Q(qn),
    .SETN(nreset)
  );
endmodule
