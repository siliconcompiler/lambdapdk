// //#############################################################################
// //# Function:  Positive edge-triggered static inverting D-type flop-flop with #
// //             async active low reset.                                        #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_dffrqn #(
//     parameter PROP = "DEFAULT"
// ) (
//     input      d,
//     input      clk,
//     input      nreset,
//     output reg qn
// );
// 
//   always @(posedge clk or negedge nreset)
//     if (!nreset) qn <= 1'b1;
//     else qn <= ~d;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_dffrqn.v:11.1-24.10" *)
module la_dffrqn (
    d,
    clk,
    nreset,
    qn
);
  (* src = "inputs/la_dffrqn.v:20.3-22.19" *)
  wire _0_;
  wire _1_;
  wire _2_;
  (* src = "inputs/la_dffrqn.v:15.16-15.19" *)
  input clk;
  wire clk;
  (* src = "inputs/la_dffrqn.v:14.16-14.17" *)
  input d;
  wire d;
  (* src = "inputs/la_dffrqn.v:16.16-16.22" *)
  input nreset;
  wire nreset;
  (* src = "inputs/la_dffrqn.v:17.16-17.18" *)
  output qn;
  wire qn;
  INVx2_ASAP7_75t_L _3_ (
      .A(d),
      .Y(_0_)
  );
  INVx2_ASAP7_75t_L _4_ (
      .A(_1_),
      .Y(qn)
  );
  (* src = "inputs/la_dffrqn.v:20.3-22.19" *)
  DFFASRHQNx1_ASAP7_75t_L _5_ (
      .CLK(clk),
      .D(_0_),
      .QN(_1_),
      .RESETN(nreset),
      .SETN(_2_)
  );
  TIEHIx1_ASAP7_75t_L _6_ (.H(_2_));
endmodule
