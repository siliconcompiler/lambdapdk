// //#############################################################################
// //# Function:  Positive edge-triggered static inverting D-type flop-flop with #
// //             async active low set.                                          #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_dffsqn #(
//     parameter PROP = "DEFAULT"
// ) (
//     input d,
//     input clk,
//     input nset,
//     output reg qn
// );
// 
//     always @(posedge clk or negedge nset)
//         if (!nset) qn <= 1'b0;
//         else qn <= ~d;
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "inputs/la_dffsqn.v:11.1-24.10" *)
module la_dffsqn (
    d,
    clk,
    nset,
    qn
);
  (* src = "inputs/la_dffsqn.v:20.5-22.23" *)
  wire _0_;
  wire _1_;
  wire _2_;
  (* src = "inputs/la_dffsqn.v:15.11-15.14" *)
  input clk;
  wire clk;
  (* src = "inputs/la_dffsqn.v:14.11-14.12" *)
  input d;
  wire d;
  (* src = "inputs/la_dffsqn.v:16.11-16.15" *)
  input nset;
  wire nset;
  (* src = "inputs/la_dffsqn.v:17.16-17.18" *)
  output qn;
  wire qn;
  INVx2_ASAP7_75t_R _3_ (
      .A(d),
      .Y(_0_)
  );
  INVx2_ASAP7_75t_R _4_ (
      .A(_1_),
      .Y(qn)
  );
  (* src = "inputs/la_dffsqn.v:20.5-22.23" *)
  DFFASRHQNx1_ASAP7_75t_R _5_ (
      .CLK(clk),
      .D(_0_),
      .QN(_1_),
      .RESETN(_2_),
      .SETN(nset)
  );
  TIEHIx1_ASAP7_75t_R _6_ (.H(_2_));
endmodule
