// //#############################################################################
// //# Function:  Reset synchronizer (async assert, sync deassert)               #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:   MIT (see LICENSE file in Lambda repository)                    #
// //#############################################################################
// 
// module la_rsync #(
//     parameter PROP = "DEFAULT"
// ) (
//     input clk,  // clock
//     input nrst_in,  // async reset input
//     output nrst_out  // async assert, sync deassert reset
// );
// 
//     localparam STAGES = 2;
//     localparam RND = 1;
// 
//     reg     [STAGES:0] sync_pipe;
//     integer            sync_delay;
// 
// `ifndef SYNTHESIS
//     always @(posedge clk) sync_delay <= {$random} % 2;
// `endif
// 
//     always @(posedge clk or negedge nrst_in)
//         if (!nrst_in) sync_pipe[STAGES:0] <= 'b0;
//         else sync_pipe[STAGES:0] <= {sync_pipe[STAGES-1:0], 1'b1};
// 
// `ifdef SYNTHESIS
//     assign nrst_out = sync_pipe[STAGES-1];
// `else
//     assign nrst_out = (|sync_delay & (|RND)) ? sync_pipe[STAGES] : sync_pipe[STAGES-1];
// `endif
// 
// endmodule

/* Generated by Yosys 0.40 (git sha1 a1bb0255d, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_rsync(clk, nrst_in, nrst_out);
  wire _0_;
  wire _1_;
  wire _2_;
  input clk;
  wire clk;
  input nrst_in;
  wire nrst_in;
  output nrst_out;
  wire nrst_out;
  wire \sync_pipe[0] ;
  INVx1_ASAP7_75t_L _3_ (
    .A(_0_),
    .Y(nrst_out)
  );
  INVx1_ASAP7_75t_L _4_ (
    .A(_1_),
    .Y(\sync_pipe[0] )
  );
  DFFASRHQNx1_ASAP7_75t_L _5_ (
    .CLK(clk),
    .D(_2_),
    .QN(_1_),
    .RESETN(_2_),
    .SETN(nrst_in)
  );
  DFFASRHQNx1_ASAP7_75t_L _6_ (
    .CLK(clk),
    .D(\sync_pipe[0] ),
    .QN(_0_),
    .RESETN(_2_),
    .SETN(nrst_in)
  );
  TIEHIx1_ASAP7_75t_L _7_ (
    .H(_2_)
  );
endmodule
