// //#############################################################################
// //# Function: Tie High Cell                                                   #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_tiehi #(
//     parameter PROP = "DEFAULT"
// ) (
//     output z
// );
// 
//     assign z = 1'b1;
// 
// endmodule

/* Generated by Yosys 0.40+33 (git sha1 cd1fb8b15, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_tiehi(z);
  output z;
  wire z;
  sg13g2_tiehi _0_ (
    .L_HI(z)
  );
endmodule
