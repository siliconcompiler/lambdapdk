// //#############################################################################
// //# Function: 2-Input Inverting Mux                                           #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_muxi2 #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  d0,
//     input  d1,
//     input  s,
//     output z
// );
// 
//     assign z = ~((d0 & ~s) | (d1 & s));
// 
// endmodule

/* Generated by Yosys 0.44 (git sha1 80ba43d26, g++ 11.4.0-1ubuntu1~22.04 -fPIC -O3) */

(* top =  1  *)
(* src = "generated" *)
module la_muxi2 (
    d0,
    d1,
    s,
    z
);
  wire _0_;
  (* src = "generated" *)
  input d0;
  wire d0;
  (* src = "generated" *)
  input d1;
  wire d1;
  (* src = "generated" *)
  input s;
  wire s;
  (* src = "generated" *)
  output z;
  wire z;
  gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1_ (
      .I0(d0),
      .I1(d1),
      .S (s),
      .Z (_0_)
  );
  gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2_ (
      .I (_0_),
      .ZN(z)
  );
endmodule
