// //#############################################################################
// //# Function: 2-Input Inverting Mux                                           #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_muxi2 #(parameter PROP = "DEFAULT")   (
//     input  d0,
//     input  d1,
//     input  s,
//     output z
//     );
// 
//    assign z = ~((d0 & ~s) | (d1 & s));
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_muxi2(d0, d1, s, z);
  wire _0_;
  input d0;
  wire d0;
  input d1;
  wire d1;
  input s;
  wire s;
  output z;
  wire z;
  gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1_ (
    .I0(d0),
    .I1(d1),
    .S(s),
    .Z(_0_)
  );
  gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2_ (
    .I(_0_),
    .ZN(z)
  );
endmodule
