// //#############################################################################
// //# Function: Synchronizer with async reset                                   #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// module la_drsync #(
//     parameter PROP = "DEFAULT"
// ) (
//     input  clk,    // clock
//     input  in,     // input data
//     input  nreset, // async active low reset
//     output out     // synchronized data
// );
// 
//     localparam STAGES = 2;
// 
//     reg [STAGES-1:0] shiftreg;
// 
//     always @(posedge clk or negedge nreset)
//         if (!nreset) shiftreg[STAGES-1:0] <= 'b0;
//         else shiftreg[STAGES-1:0] <= {shiftreg[STAGES-2:0], in};
// 
//     assign out = shiftreg[STAGES-1];
// 
// endmodule

/* Generated by Yosys 0.40 (git sha1 a1bb0255d, g++ 11.4.0-1ubuntu1~22.04 -fPIC -Os) */

module la_drsync(clk, in, nreset, out);
  wire _0_;
  wire _1_;
  wire _2_;
  input clk;
  wire clk;
  input in;
  wire in;
  input nreset;
  wire nreset;
  output out;
  wire out;
  wire \shiftreg[0] ;
  INVx1_ASAP7_75t_SL _3_ (
    .A(_0_),
    .Y(out)
  );
  INVx1_ASAP7_75t_SL _4_ (
    .A(_1_),
    .Y(\shiftreg[0] )
  );
  DFFASRHQNx1_ASAP7_75t_SL _5_ (
    .CLK(clk),
    .D(in),
    .QN(_1_),
    .RESETN(_2_),
    .SETN(nreset)
  );
  DFFASRHQNx1_ASAP7_75t_SL _6_ (
    .CLK(clk),
    .D(\shiftreg[0] ),
    .QN(_0_),
    .RESETN(_2_),
    .SETN(nreset)
  );
  TIEHIx1_ASAP7_75t_SL _7_ (
    .H(_2_)
  );
endmodule
