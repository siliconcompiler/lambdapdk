// //#############################################################################
// //# Function: Integrated "And" Clock Gating Cell (And)                        #
// //# Copyright: Lambda Project Authors. All rights Reserved.                   #
// //# License:  MIT (see LICENSE file in Lambda repository)                     #
// //#############################################################################
// 
// module la_clkicgand #(parameter PROP = "DEFAULT")  (
//    input  clk, // clock input
//    input  te, // test enable
//    input  en, // enable (from positive edge FF)
//    output eclk // enabled clock output
//    );
// 
//    reg 	  en_stable;
// 
//    always @ (clk or en or te)
//      if (~clk)
//        en_stable <= en | te;
// 
//    assign eclk =  clk & en_stable;
// 
// endmodule

/* Generated by Yosys 0.37 (git sha1 a5c7f69ed, clang 14.0.0-1ubuntu1.1 -fPIC -Os) */

module la_clkicgand(clk, te, en, eclk);
  wire _0_;
  wire _1_;
  input clk;
  wire clk;
  output eclk;
  wire eclk;
  input en;
  wire en;
  wire en_stable;
  input te;
  wire te;
  gf180mcu_fd_sc_mcu9t5v0__and2_2 _2_ (
    .A1(en_stable),
    .A2(clk),
    .Z(eclk)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_2 _3_ (
    .A1(te),
    .A2(en),
    .Z(_0_)
  );
  gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _4_ (
    .I(clk),
    .ZN(_1_)
  );
  gf180mcu_fd_sc_mcu9t5v0__latq_1 _5_ (
    .D(_0_),
    .E(_1_),
    .Q(en_stable)
  );
endmodule
